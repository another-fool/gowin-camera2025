module gw_gao(
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[27] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[26] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[25] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[24] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[23] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[22] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[21] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[20] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[19] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[18] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[17] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[16] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[15] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[14] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[13] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[12] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[11] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[10] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[9] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[8] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[7] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[6] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[5] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[4] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[3] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[2] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[1] ,
    \mux_top_inst/algorithm_top_inst/current_buffer_addr[0] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[28] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[27] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[26] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[25] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[24] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[23] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[22] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[21] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[20] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[19] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[18] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[17] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[16] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[15] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[14] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[13] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[12] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[11] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[10] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[9] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[8] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[7] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[6] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[5] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[4] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[3] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[2] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[1] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[0] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[15] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[14] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[13] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[12] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[11] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[10] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[9] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[8] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[7] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[6] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[5] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[4] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[3] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[2] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[1] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[0] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[255] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[254] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[253] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[252] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[251] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[250] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[249] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[248] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[247] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[246] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[245] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[244] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[243] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[242] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[241] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[240] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[239] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[238] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[237] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[236] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[235] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[234] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[233] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[232] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[231] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[230] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[229] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[228] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[227] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[226] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[225] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[224] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[223] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[222] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[221] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[220] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[219] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[218] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[217] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[216] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[215] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[214] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[213] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[212] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[211] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[210] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[209] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[208] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[207] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[206] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[205] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[204] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[203] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[202] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[201] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[200] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[199] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[198] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[197] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[196] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[195] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[194] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[193] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[192] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[191] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[190] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[189] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[188] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[187] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[186] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[185] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[184] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[183] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[182] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[181] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[180] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[179] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[178] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[177] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[176] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[175] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[174] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[173] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[172] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[171] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[170] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[169] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[168] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[167] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[166] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[165] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[164] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[163] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[162] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[161] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[160] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[159] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[158] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[157] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[156] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[155] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[154] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[153] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[152] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[151] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[150] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[149] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[148] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[147] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[146] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[145] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[144] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[143] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[142] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[141] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[140] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[139] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[138] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[137] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[136] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[135] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[134] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[133] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[132] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[131] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[130] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[129] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[128] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[127] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[126] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[125] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[124] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[123] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[122] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[121] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[120] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[119] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[118] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[117] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[116] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[115] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[114] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[113] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[112] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[111] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[110] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[109] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[108] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[107] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[106] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[105] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[104] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[103] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[102] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[101] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[100] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[99] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[98] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[97] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[96] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[95] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[94] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[93] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[92] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[91] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[90] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[89] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[88] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[87] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[86] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[85] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[84] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[83] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[82] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[81] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[80] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[79] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[78] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[77] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[76] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[75] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[74] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[73] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[72] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[71] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[70] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[69] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[68] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[67] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[66] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[65] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[64] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[63] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[62] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[61] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[60] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[59] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[58] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[57] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[56] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[55] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[54] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[53] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[52] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[51] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[50] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[49] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[48] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[47] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[46] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[45] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[44] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[43] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[42] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[41] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[40] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[39] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[38] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[37] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[36] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[35] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[34] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[33] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[32] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[31] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[30] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[29] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[28] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[27] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[26] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[25] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[24] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[23] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[22] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[21] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[20] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[19] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[18] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[17] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[16] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[15] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[14] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[13] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[12] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[11] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[10] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[9] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[8] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[7] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[6] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[5] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[4] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[3] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[2] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[1] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[0] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[28] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[27] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[26] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[25] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[24] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[23] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[22] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[21] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[20] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[19] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[18] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[17] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[16] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[15] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[14] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[13] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[12] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[11] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[10] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[9] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[8] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[7] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[6] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[5] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[4] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[3] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[2] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[1] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[0] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[15] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[14] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[13] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[12] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[11] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[10] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[9] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[8] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[7] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[6] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[5] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[4] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[3] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[2] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[1] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[0] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[255] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[254] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[253] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[252] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[251] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[250] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[249] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[248] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[247] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[246] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[245] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[244] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[243] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[242] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[241] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[240] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[239] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[238] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[237] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[236] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[235] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[234] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[233] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[232] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[231] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[230] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[229] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[228] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[227] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[226] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[225] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[224] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[223] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[222] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[221] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[220] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[219] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[218] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[217] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[216] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[215] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[214] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[213] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[212] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[211] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[210] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[209] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[208] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[207] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[206] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[205] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[204] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[203] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[202] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[201] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[200] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[199] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[198] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[197] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[196] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[195] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[194] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[193] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[192] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[191] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[190] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[189] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[188] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[187] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[186] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[185] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[184] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[183] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[182] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[181] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[180] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[179] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[178] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[177] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[176] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[175] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[174] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[173] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[172] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[171] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[170] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[169] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[168] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[167] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[166] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[165] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[164] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[163] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[162] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[161] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[160] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[159] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[158] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[157] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[156] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[155] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[154] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[153] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[152] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[151] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[150] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[149] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[148] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[147] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[146] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[145] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[144] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[143] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[142] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[141] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[140] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[139] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[138] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[137] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[136] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[135] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[134] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[133] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[132] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[131] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[130] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[129] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[128] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[127] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[126] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[125] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[124] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[123] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[122] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[121] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[120] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[119] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[118] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[117] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[116] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[115] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[114] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[113] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[112] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[111] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[110] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[109] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[108] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[107] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[106] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[105] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[104] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[103] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[102] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[101] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[100] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[99] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[98] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[97] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[96] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[95] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[94] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[93] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[92] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[91] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[90] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[89] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[88] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[87] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[86] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[85] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[84] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[83] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[82] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[81] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[80] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[79] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[78] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[77] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[76] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[75] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[74] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[73] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[72] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[71] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[70] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[69] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[68] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[67] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[66] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[65] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[64] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[63] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[62] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[61] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[60] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[59] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[58] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[57] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[56] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[55] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[54] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[53] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[52] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[51] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[50] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[49] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[48] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[47] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[46] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[45] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[44] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[43] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[42] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[41] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[40] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[39] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[38] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[37] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[36] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[35] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[34] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[33] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[32] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[31] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[30] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[29] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[28] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[27] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[26] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[25] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[24] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[23] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[22] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[21] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[20] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[19] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[18] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[17] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[16] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[15] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[14] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[13] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[12] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[11] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[10] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[9] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[8] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[7] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[6] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[5] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[4] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[3] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[2] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[1] ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[0] ,
    \mux_top_inst/algorithm_top_inst/time_out[19] ,
    \mux_top_inst/algorithm_top_inst/time_out[18] ,
    \mux_top_inst/algorithm_top_inst/time_out[17] ,
    \mux_top_inst/algorithm_top_inst/time_out[16] ,
    \mux_top_inst/algorithm_top_inst/time_out[15] ,
    \mux_top_inst/algorithm_top_inst/time_out[14] ,
    \mux_top_inst/algorithm_top_inst/time_out[13] ,
    \mux_top_inst/algorithm_top_inst/time_out[12] ,
    \mux_top_inst/algorithm_top_inst/time_out[11] ,
    \mux_top_inst/algorithm_top_inst/time_out[10] ,
    \mux_top_inst/algorithm_top_inst/time_out[9] ,
    \mux_top_inst/algorithm_top_inst/time_out[8] ,
    \mux_top_inst/algorithm_top_inst/time_out[7] ,
    \mux_top_inst/algorithm_top_inst/time_out[6] ,
    \mux_top_inst/algorithm_top_inst/time_out[5] ,
    \mux_top_inst/algorithm_top_inst/time_out[4] ,
    \mux_top_inst/algorithm_top_inst/time_out[3] ,
    \mux_top_inst/algorithm_top_inst/time_out[2] ,
    \mux_top_inst/algorithm_top_inst/time_out[1] ,
    \mux_top_inst/algorithm_top_inst/time_out[0] ,
    \mux_top_inst/algorithm_top_inst/cs[7] ,
    \mux_top_inst/algorithm_top_inst/cs[6] ,
    \mux_top_inst/algorithm_top_inst/cs[5] ,
    \mux_top_inst/algorithm_top_inst/cs[4] ,
    \mux_top_inst/algorithm_top_inst/cs[3] ,
    \mux_top_inst/algorithm_top_inst/cs[2] ,
    \mux_top_inst/algorithm_top_inst/cs[1] ,
    \mux_top_inst/algorithm_top_inst/cs[0] ,
    \mux_top_inst/algorithm_top_inst/cmos_cnt[4] ,
    \mux_top_inst/algorithm_top_inst/cmos_cnt[3] ,
    \mux_top_inst/algorithm_top_inst/cmos_cnt[2] ,
    \mux_top_inst/algorithm_top_inst/cmos_cnt[1] ,
    \mux_top_inst/algorithm_top_inst/cmos_cnt[0] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[10] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[9] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[8] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[7] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[6] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[5] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[4] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[3] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[2] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[1] ,
    \mux_top_inst/algorithm_top_inst/line_cnt[0] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[255] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[254] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[253] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[252] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[251] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[250] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[249] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[248] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[247] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[246] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[245] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[244] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[243] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[242] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[241] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[240] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[239] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[238] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[237] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[236] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[235] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[234] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[233] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[232] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[231] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[230] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[229] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[228] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[227] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[226] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[225] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[224] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[223] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[222] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[221] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[220] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[219] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[218] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[217] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[216] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[215] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[214] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[213] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[212] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[211] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[210] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[209] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[208] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[207] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[206] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[205] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[204] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[203] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[202] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[201] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[200] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[199] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[198] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[197] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[196] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[195] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[194] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[193] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[192] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[191] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[190] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[189] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[188] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[187] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[186] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[185] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[184] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[183] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[182] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[181] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[180] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[179] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[178] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[177] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[176] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[175] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[174] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[173] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[172] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[171] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[170] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[169] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[168] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[167] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[166] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[165] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[164] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[163] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[162] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[161] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[160] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[159] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[158] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[157] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[156] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[155] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[154] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[153] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[152] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[151] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[150] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[149] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[148] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[147] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[146] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[145] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[144] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[143] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[142] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[141] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[140] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[139] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[138] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[137] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[136] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[135] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[134] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[133] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[132] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[131] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[130] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[129] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[128] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[127] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[126] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[125] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[124] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[123] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[122] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[121] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[120] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[119] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[118] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[117] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[116] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[115] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[114] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[113] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[112] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[111] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[110] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[109] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[108] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[107] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[106] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[105] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[104] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[103] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[102] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[101] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[100] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[99] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[98] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[97] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[96] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[95] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[94] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[93] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[92] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[91] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[90] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[89] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[88] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[87] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[86] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[85] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[84] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[83] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[82] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[81] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[80] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[79] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[78] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[77] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[76] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[75] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[74] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[73] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[72] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[71] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[70] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[69] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[68] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[67] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[66] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[65] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[64] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[63] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[62] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[61] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[60] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[59] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[58] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[57] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[56] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[55] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[54] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[53] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[52] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[51] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[50] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[49] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[48] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[47] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[46] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[45] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[44] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[43] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[42] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[41] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[40] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[39] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[38] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[37] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[36] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[35] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[34] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[33] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[32] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[31] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[30] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[29] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[28] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[27] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[26] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[25] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[24] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[23] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[22] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[21] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[20] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[19] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[18] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[17] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[16] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[15] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[14] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[13] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[12] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[11] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[10] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[9] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[8] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[7] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[6] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[5] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[4] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[3] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[2] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[1] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_data[0] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[255] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[254] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[253] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[252] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[251] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[250] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[249] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[248] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[247] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[246] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[245] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[244] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[243] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[242] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[241] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[240] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[239] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[238] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[237] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[236] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[235] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[234] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[233] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[232] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[231] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[230] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[229] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[228] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[227] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[226] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[225] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[224] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[223] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[222] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[221] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[220] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[219] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[218] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[217] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[216] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[215] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[214] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[213] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[212] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[211] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[210] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[209] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[208] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[207] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[206] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[205] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[204] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[203] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[202] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[201] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[200] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[199] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[198] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[197] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[196] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[195] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[194] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[193] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[192] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[191] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[190] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[189] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[188] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[187] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[186] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[185] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[184] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[183] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[182] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[181] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[180] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[179] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[178] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[177] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[176] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[175] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[174] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[173] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[172] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[171] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[170] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[169] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[168] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[167] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[166] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[165] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[164] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[163] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[162] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[161] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[160] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[159] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[158] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[157] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[156] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[155] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[154] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[153] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[152] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[151] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[150] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[149] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[148] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[147] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[146] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[145] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[144] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[143] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[142] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[141] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[140] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[139] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[138] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[137] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[136] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[135] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[134] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[133] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[132] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[131] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[130] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[129] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[128] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[127] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[126] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[125] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[124] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[123] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[122] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[121] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[120] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[119] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[118] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[117] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[116] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[115] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[114] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[113] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[112] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[111] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[110] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[109] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[108] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[107] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[106] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[105] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[104] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[103] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[102] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[101] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[100] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[99] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[98] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[97] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[96] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[95] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[94] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[93] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[92] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[91] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[90] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[89] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[88] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[87] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[86] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[85] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[84] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[83] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[82] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[81] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[80] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[79] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[78] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[77] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[76] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[75] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[74] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[73] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[72] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[71] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[70] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[69] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[68] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[67] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[66] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[65] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[64] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[63] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[62] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[61] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[60] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[59] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[58] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[57] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[56] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[55] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[54] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[53] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[52] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[51] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[50] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[49] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[48] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[47] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[46] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[45] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[44] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[43] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[42] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[41] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[40] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[39] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[38] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[37] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[36] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[35] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[34] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[33] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[32] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[31] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[30] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[29] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[28] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[27] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[26] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[25] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[24] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[23] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[22] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[21] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[20] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[19] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[18] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[17] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[16] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[15] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[14] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[13] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[12] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[11] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[10] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[9] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[8] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[7] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[6] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[5] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[4] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[3] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[2] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[1] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_data[0] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[6] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[5] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[4] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[3] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[2] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[1] ,
    \mux_top_inst/algorithm_top_inst/ram_wr_addr[0] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[6] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[5] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[4] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[3] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[2] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[1] ,
    \mux_top_inst/algorithm_top_inst/ram_rd_addr[0] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[27] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[26] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[25] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[24] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[23] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[22] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[21] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[20] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[19] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[18] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[17] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[16] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[15] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[14] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[13] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[12] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[11] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[10] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[9] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[8] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[7] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[6] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[5] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[4] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[3] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[2] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[1] ,
    \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[0] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[27] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[26] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[25] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[24] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[23] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[22] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[21] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[20] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[19] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[18] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[17] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[16] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[15] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[14] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[13] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[12] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[11] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[10] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[9] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[8] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[7] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[6] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[5] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[4] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[3] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[2] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[1] ,
    \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[0] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[27] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[26] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[25] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[24] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[23] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[22] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[21] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[20] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[19] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[18] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[17] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[16] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[15] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[14] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[13] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[12] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[11] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[10] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[9] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[8] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[7] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[6] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[5] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[4] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[3] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[2] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[1] ,
    \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[0] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[11] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[10] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[9] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[8] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[7] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[6] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[5] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[4] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[3] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[2] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[1] ,
    \mux_top_inst/algorithm_top_inst/cnt_rx_pix[0] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[27] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[26] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[25] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[24] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[23] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[22] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[21] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[20] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[19] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[18] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[17] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[16] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[15] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[14] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[13] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[12] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[11] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[10] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[9] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[8] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[7] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[6] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[5] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[4] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[3] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[2] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[1] ,
    \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[0] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[255] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[254] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[253] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[252] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[251] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[250] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[249] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[248] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[247] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[246] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[245] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[244] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[243] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[242] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[241] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[240] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[239] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[238] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[237] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[236] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[235] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[234] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[233] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[232] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[231] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[230] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[229] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[228] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[227] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[226] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[225] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[224] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[223] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[222] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[221] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[220] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[219] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[218] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[217] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[216] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[215] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[214] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[213] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[212] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[211] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[210] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[209] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[208] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[207] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[206] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[205] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[204] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[203] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[202] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[201] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[200] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[199] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[198] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[197] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[196] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[195] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[194] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[193] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[192] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[191] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[190] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[189] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[188] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[187] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[186] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[185] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[184] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[183] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[182] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[181] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[180] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[179] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[178] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[177] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[176] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[175] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[174] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[173] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[172] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[171] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[170] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[169] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[168] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[167] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[166] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[165] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[164] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[163] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[162] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[161] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[160] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[159] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[158] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[157] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[156] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[155] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[154] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[153] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[152] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[151] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[150] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[149] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[148] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[147] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[146] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[145] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[144] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[143] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[142] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[141] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[140] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[139] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[138] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[137] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[136] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[135] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[134] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[133] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[132] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[131] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[130] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[129] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[128] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[127] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[126] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[125] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[124] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[123] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[122] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[121] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[120] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[119] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[118] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[117] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[116] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[115] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[114] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[113] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[112] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[111] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[110] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[109] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[108] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[107] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[106] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[105] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[104] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[103] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[102] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[101] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[100] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[99] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[98] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[97] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[96] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[95] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[94] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[93] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[92] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[91] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[90] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[89] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[88] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[87] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[86] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[85] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[84] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[83] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[82] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[81] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[80] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[79] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[78] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[77] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[76] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[75] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[74] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[73] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[72] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[71] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[70] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[69] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[68] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[67] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[66] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[65] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[64] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[63] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[62] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[61] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[60] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[59] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[58] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[57] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[56] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[55] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[54] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[53] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[52] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[51] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[50] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[49] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[48] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[47] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[46] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[45] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[44] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[43] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[42] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[41] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[40] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[39] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[38] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[37] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[36] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[35] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[34] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[33] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[32] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[31] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[30] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[29] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[28] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[27] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[26] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[25] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[24] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[23] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[22] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[21] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[20] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[19] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[18] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[17] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[16] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[15] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[14] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[13] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[12] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[11] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[10] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[9] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[8] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[7] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[6] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[5] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[4] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[3] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[2] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[1] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/dout[0] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[6] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[5] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[4] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[3] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[2] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[1] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ada[0] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[255] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[254] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[253] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[252] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[251] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[250] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[249] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[248] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[247] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[246] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[245] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[244] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[243] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[242] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[241] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[240] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[239] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[238] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[237] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[236] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[235] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[234] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[233] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[232] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[231] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[230] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[229] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[228] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[227] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[226] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[225] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[224] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[223] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[222] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[221] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[220] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[219] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[218] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[217] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[216] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[215] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[214] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[213] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[212] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[211] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[210] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[209] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[208] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[207] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[206] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[205] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[204] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[203] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[202] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[201] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[200] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[199] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[198] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[197] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[196] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[195] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[194] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[193] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[192] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[191] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[190] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[189] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[188] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[187] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[186] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[185] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[184] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[183] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[182] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[181] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[180] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[179] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[178] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[177] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[176] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[175] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[174] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[173] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[172] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[171] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[170] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[169] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[168] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[167] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[166] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[165] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[164] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[163] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[162] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[161] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[160] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[159] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[158] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[157] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[156] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[155] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[154] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[153] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[152] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[151] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[150] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[149] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[148] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[147] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[146] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[145] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[144] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[143] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[142] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[141] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[140] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[139] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[138] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[137] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[136] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[135] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[134] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[133] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[132] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[131] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[130] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[129] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[128] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[127] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[126] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[125] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[124] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[123] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[122] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[121] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[120] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[119] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[118] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[117] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[116] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[115] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[114] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[113] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[112] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[111] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[110] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[109] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[108] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[107] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[106] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[105] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[104] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[103] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[102] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[101] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[100] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[99] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[98] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[97] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[96] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[95] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[94] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[93] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[92] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[91] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[90] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[89] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[88] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[87] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[86] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[85] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[84] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[83] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[82] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[81] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[80] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[79] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[78] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[77] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[76] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[75] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[74] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[73] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[72] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[71] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[70] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[69] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[68] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[67] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[66] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[65] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[64] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[63] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[62] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[61] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[60] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[59] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[58] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[57] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[56] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[55] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[54] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[53] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[52] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[51] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[50] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[49] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[48] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[47] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[46] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[45] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[44] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[43] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[42] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[41] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[40] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[39] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[38] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[37] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[36] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[35] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[34] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[33] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[32] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[31] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[30] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[29] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[28] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[27] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[26] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[25] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[24] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[23] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[22] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[21] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[20] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[19] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[18] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[17] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[16] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[15] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[14] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[13] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[12] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[11] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[10] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[9] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[8] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[7] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[6] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[5] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[4] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[3] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[2] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[1] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/din[0] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[6] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[5] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[4] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[3] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[2] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[1] ,
    \mux_top_inst/algorithm_top_inst/buffer_line/adb[0] ,
    \mux_top_inst/algorithm_top_inst/syn_off0_vs ,
    \mux_top_inst/algorithm_top_inst/coms0_wr_area ,
    \mux_top_inst/algorithm_top_inst/coms1_wr_area ,
    \mux_top_inst/algorithm_top_inst/coms2_wr_area ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.req ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.finish ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.ack ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.data_req ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.req ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.ack ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.dv ,
    \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.finish ,
    \mux_top_inst/algorithm_top_inst/cs_r1 ,
    \mux_top_inst/algorithm_top_inst/cs_r2 ,
    \mux_top_inst/algorithm_top_inst/cs_rise ,
    \mux_top_inst/algorithm_top_inst/ram_rd_en ,
    \mux_top_inst/algorithm_top_inst/ram_wr_en ,
    \mux_top_inst/algorithm_top_inst/buffer_line/clka ,
    \mux_top_inst/algorithm_top_inst/buffer_line/cea ,
    \mux_top_inst/algorithm_top_inst/buffer_line/clkb ,
    \mux_top_inst/algorithm_top_inst/buffer_line/ceb ,
    \mux_top_inst/algorithm_top_inst/buffer_line/oce ,
    \mux_top_inst/algorithm_top_inst/buffer_line/reset ,
    \mux_top_inst/hdmi_rd_inst/ddr_clk ,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \mux_top_inst/algorithm_top_inst/current_buffer_addr[27] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[26] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[25] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[24] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[23] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[22] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[21] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[20] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[19] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[18] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[17] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[16] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[15] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[14] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[13] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[12] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[11] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[10] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[9] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[8] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[7] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[6] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[5] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[4] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[3] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[2] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[1] ;
input \mux_top_inst/algorithm_top_inst/current_buffer_addr[0] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[28] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[27] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[26] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[25] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[24] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[23] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[22] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[21] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[20] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[19] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[18] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[17] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[16] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[15] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[14] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[13] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[12] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[11] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[10] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[9] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[8] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[7] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[6] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[5] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[4] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[3] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[2] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[1] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[0] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[15] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[14] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[13] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[12] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[11] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[10] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[9] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[8] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[7] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[6] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[5] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[4] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[3] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[2] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[1] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[0] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[255] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[254] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[253] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[252] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[251] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[250] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[249] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[248] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[247] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[246] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[245] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[244] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[243] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[242] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[241] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[240] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[239] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[238] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[237] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[236] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[235] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[234] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[233] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[232] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[231] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[230] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[229] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[228] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[227] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[226] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[225] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[224] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[223] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[222] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[221] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[220] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[219] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[218] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[217] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[216] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[215] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[214] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[213] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[212] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[211] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[210] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[209] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[208] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[207] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[206] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[205] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[204] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[203] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[202] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[201] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[200] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[199] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[198] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[197] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[196] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[195] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[194] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[193] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[192] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[191] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[190] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[189] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[188] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[187] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[186] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[185] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[184] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[183] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[182] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[181] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[180] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[179] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[178] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[177] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[176] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[175] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[174] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[173] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[172] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[171] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[170] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[169] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[168] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[167] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[166] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[165] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[164] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[163] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[162] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[161] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[160] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[159] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[158] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[157] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[156] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[155] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[154] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[153] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[152] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[151] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[150] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[149] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[148] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[147] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[146] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[145] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[144] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[143] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[142] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[141] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[140] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[139] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[138] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[137] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[136] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[135] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[134] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[133] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[132] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[131] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[130] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[129] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[128] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[127] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[126] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[125] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[124] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[123] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[122] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[121] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[120] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[119] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[118] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[117] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[116] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[115] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[114] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[113] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[112] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[111] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[110] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[109] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[108] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[107] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[106] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[105] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[104] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[103] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[102] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[101] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[100] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[99] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[98] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[97] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[96] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[95] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[94] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[93] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[92] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[91] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[90] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[89] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[88] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[87] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[86] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[85] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[84] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[83] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[82] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[81] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[80] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[79] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[78] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[77] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[76] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[75] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[74] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[73] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[72] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[71] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[70] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[69] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[68] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[67] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[66] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[65] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[64] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[63] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[62] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[61] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[60] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[59] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[58] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[57] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[56] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[55] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[54] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[53] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[52] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[51] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[50] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[49] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[48] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[47] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[46] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[45] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[44] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[43] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[42] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[41] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[40] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[39] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[38] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[37] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[36] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[35] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[34] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[33] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[32] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[31] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[30] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[29] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[28] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[27] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[26] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[25] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[24] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[23] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[22] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[21] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[20] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[19] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[18] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[17] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[16] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[15] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[14] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[13] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[12] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[11] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[10] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[9] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[8] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[7] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[6] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[5] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[4] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[3] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[2] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[1] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[0] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[28] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[27] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[26] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[25] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[24] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[23] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[22] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[21] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[20] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[19] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[18] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[17] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[16] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[15] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[14] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[13] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[12] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[11] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[10] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[9] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[8] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[7] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[6] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[5] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[4] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[3] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[2] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[1] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[0] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[15] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[14] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[13] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[12] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[11] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[10] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[9] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[8] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[7] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[6] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[5] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[4] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[3] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[2] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[1] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[0] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[255] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[254] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[253] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[252] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[251] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[250] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[249] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[248] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[247] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[246] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[245] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[244] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[243] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[242] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[241] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[240] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[239] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[238] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[237] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[236] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[235] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[234] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[233] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[232] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[231] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[230] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[229] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[228] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[227] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[226] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[225] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[224] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[223] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[222] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[221] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[220] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[219] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[218] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[217] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[216] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[215] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[214] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[213] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[212] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[211] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[210] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[209] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[208] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[207] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[206] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[205] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[204] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[203] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[202] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[201] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[200] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[199] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[198] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[197] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[196] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[195] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[194] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[193] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[192] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[191] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[190] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[189] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[188] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[187] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[186] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[185] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[184] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[183] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[182] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[181] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[180] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[179] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[178] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[177] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[176] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[175] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[174] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[173] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[172] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[171] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[170] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[169] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[168] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[167] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[166] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[165] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[164] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[163] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[162] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[161] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[160] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[159] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[158] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[157] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[156] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[155] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[154] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[153] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[152] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[151] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[150] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[149] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[148] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[147] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[146] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[145] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[144] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[143] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[142] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[141] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[140] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[139] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[138] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[137] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[136] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[135] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[134] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[133] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[132] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[131] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[130] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[129] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[128] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[127] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[126] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[125] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[124] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[123] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[122] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[121] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[120] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[119] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[118] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[117] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[116] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[115] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[114] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[113] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[112] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[111] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[110] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[109] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[108] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[107] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[106] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[105] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[104] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[103] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[102] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[101] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[100] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[99] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[98] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[97] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[96] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[95] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[94] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[93] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[92] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[91] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[90] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[89] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[88] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[87] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[86] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[85] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[84] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[83] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[82] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[81] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[80] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[79] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[78] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[77] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[76] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[75] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[74] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[73] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[72] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[71] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[70] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[69] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[68] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[67] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[66] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[65] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[64] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[63] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[62] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[61] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[60] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[59] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[58] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[57] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[56] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[55] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[54] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[53] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[52] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[51] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[50] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[49] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[48] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[47] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[46] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[45] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[44] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[43] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[42] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[41] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[40] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[39] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[38] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[37] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[36] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[35] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[34] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[33] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[32] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[31] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[30] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[29] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[28] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[27] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[26] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[25] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[24] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[23] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[22] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[21] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[20] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[19] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[18] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[17] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[16] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[15] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[14] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[13] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[12] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[11] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[10] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[9] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[8] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[7] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[6] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[5] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[4] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[3] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[2] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[1] ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[0] ;
input \mux_top_inst/algorithm_top_inst/time_out[19] ;
input \mux_top_inst/algorithm_top_inst/time_out[18] ;
input \mux_top_inst/algorithm_top_inst/time_out[17] ;
input \mux_top_inst/algorithm_top_inst/time_out[16] ;
input \mux_top_inst/algorithm_top_inst/time_out[15] ;
input \mux_top_inst/algorithm_top_inst/time_out[14] ;
input \mux_top_inst/algorithm_top_inst/time_out[13] ;
input \mux_top_inst/algorithm_top_inst/time_out[12] ;
input \mux_top_inst/algorithm_top_inst/time_out[11] ;
input \mux_top_inst/algorithm_top_inst/time_out[10] ;
input \mux_top_inst/algorithm_top_inst/time_out[9] ;
input \mux_top_inst/algorithm_top_inst/time_out[8] ;
input \mux_top_inst/algorithm_top_inst/time_out[7] ;
input \mux_top_inst/algorithm_top_inst/time_out[6] ;
input \mux_top_inst/algorithm_top_inst/time_out[5] ;
input \mux_top_inst/algorithm_top_inst/time_out[4] ;
input \mux_top_inst/algorithm_top_inst/time_out[3] ;
input \mux_top_inst/algorithm_top_inst/time_out[2] ;
input \mux_top_inst/algorithm_top_inst/time_out[1] ;
input \mux_top_inst/algorithm_top_inst/time_out[0] ;
input \mux_top_inst/algorithm_top_inst/cs[7] ;
input \mux_top_inst/algorithm_top_inst/cs[6] ;
input \mux_top_inst/algorithm_top_inst/cs[5] ;
input \mux_top_inst/algorithm_top_inst/cs[4] ;
input \mux_top_inst/algorithm_top_inst/cs[3] ;
input \mux_top_inst/algorithm_top_inst/cs[2] ;
input \mux_top_inst/algorithm_top_inst/cs[1] ;
input \mux_top_inst/algorithm_top_inst/cs[0] ;
input \mux_top_inst/algorithm_top_inst/cmos_cnt[4] ;
input \mux_top_inst/algorithm_top_inst/cmos_cnt[3] ;
input \mux_top_inst/algorithm_top_inst/cmos_cnt[2] ;
input \mux_top_inst/algorithm_top_inst/cmos_cnt[1] ;
input \mux_top_inst/algorithm_top_inst/cmos_cnt[0] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[10] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[9] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[8] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[7] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[6] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[5] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[4] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[3] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[2] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[1] ;
input \mux_top_inst/algorithm_top_inst/line_cnt[0] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[255] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[254] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[253] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[252] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[251] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[250] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[249] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[248] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[247] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[246] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[245] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[244] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[243] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[242] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[241] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[240] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[239] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[238] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[237] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[236] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[235] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[234] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[233] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[232] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[231] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[230] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[229] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[228] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[227] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[226] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[225] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[224] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[223] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[222] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[221] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[220] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[219] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[218] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[217] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[216] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[215] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[214] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[213] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[212] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[211] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[210] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[209] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[208] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[207] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[206] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[205] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[204] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[203] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[202] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[201] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[200] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[199] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[198] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[197] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[196] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[195] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[194] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[193] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[192] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[191] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[190] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[189] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[188] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[187] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[186] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[185] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[184] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[183] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[182] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[181] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[180] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[179] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[178] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[177] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[176] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[175] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[174] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[173] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[172] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[171] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[170] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[169] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[168] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[167] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[166] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[165] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[164] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[163] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[162] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[161] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[160] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[159] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[158] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[157] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[156] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[155] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[154] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[153] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[152] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[151] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[150] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[149] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[148] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[147] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[146] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[145] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[144] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[143] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[142] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[141] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[140] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[139] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[138] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[137] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[136] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[135] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[134] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[133] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[132] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[131] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[130] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[129] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[128] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[127] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[126] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[125] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[124] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[123] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[122] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[121] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[120] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[119] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[118] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[117] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[116] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[115] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[114] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[113] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[112] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[111] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[110] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[109] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[108] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[107] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[106] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[105] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[104] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[103] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[102] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[101] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[100] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[99] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[98] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[97] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[96] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[95] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[94] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[93] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[92] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[91] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[90] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[89] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[88] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[87] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[86] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[85] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[84] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[83] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[82] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[81] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[80] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[79] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[78] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[77] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[76] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[75] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[74] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[73] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[72] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[71] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[70] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[69] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[68] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[67] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[66] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[65] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[64] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[63] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[62] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[61] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[60] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[59] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[58] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[57] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[56] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[55] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[54] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[53] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[52] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[51] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[50] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[49] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[48] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[47] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[46] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[45] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[44] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[43] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[42] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[41] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[40] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[39] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[38] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[37] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[36] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[35] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[34] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[33] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[32] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[31] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[30] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[29] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[28] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[27] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[26] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[25] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[24] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[23] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[22] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[21] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[20] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[19] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[18] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[17] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[16] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[15] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[14] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[13] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[12] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[11] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[10] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[9] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[8] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[7] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[6] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[5] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[4] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[3] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[2] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[1] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_data[0] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[255] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[254] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[253] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[252] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[251] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[250] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[249] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[248] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[247] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[246] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[245] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[244] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[243] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[242] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[241] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[240] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[239] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[238] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[237] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[236] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[235] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[234] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[233] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[232] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[231] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[230] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[229] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[228] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[227] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[226] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[225] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[224] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[223] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[222] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[221] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[220] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[219] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[218] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[217] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[216] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[215] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[214] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[213] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[212] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[211] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[210] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[209] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[208] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[207] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[206] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[205] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[204] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[203] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[202] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[201] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[200] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[199] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[198] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[197] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[196] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[195] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[194] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[193] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[192] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[191] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[190] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[189] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[188] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[187] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[186] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[185] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[184] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[183] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[182] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[181] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[180] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[179] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[178] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[177] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[176] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[175] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[174] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[173] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[172] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[171] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[170] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[169] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[168] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[167] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[166] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[165] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[164] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[163] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[162] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[161] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[160] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[159] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[158] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[157] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[156] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[155] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[154] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[153] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[152] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[151] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[150] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[149] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[148] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[147] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[146] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[145] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[144] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[143] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[142] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[141] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[140] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[139] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[138] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[137] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[136] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[135] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[134] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[133] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[132] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[131] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[130] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[129] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[128] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[127] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[126] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[125] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[124] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[123] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[122] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[121] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[120] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[119] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[118] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[117] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[116] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[115] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[114] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[113] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[112] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[111] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[110] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[109] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[108] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[107] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[106] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[105] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[104] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[103] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[102] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[101] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[100] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[99] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[98] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[97] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[96] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[95] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[94] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[93] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[92] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[91] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[90] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[89] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[88] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[87] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[86] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[85] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[84] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[83] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[82] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[81] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[80] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[79] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[78] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[77] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[76] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[75] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[74] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[73] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[72] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[71] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[70] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[69] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[68] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[67] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[66] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[65] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[64] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[63] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[62] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[61] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[60] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[59] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[58] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[57] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[56] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[55] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[54] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[53] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[52] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[51] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[50] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[49] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[48] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[47] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[46] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[45] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[44] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[43] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[42] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[41] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[40] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[39] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[38] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[37] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[36] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[35] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[34] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[33] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[32] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[31] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[30] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[29] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[28] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[27] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[26] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[25] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[24] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[23] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[22] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[21] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[20] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[19] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[18] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[17] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[16] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[15] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[14] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[13] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[12] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[11] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[10] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[9] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[8] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[7] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[6] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[5] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[4] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[3] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[2] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[1] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_data[0] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[6] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[5] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[4] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[3] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[2] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[1] ;
input \mux_top_inst/algorithm_top_inst/ram_wr_addr[0] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[6] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[5] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[4] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[3] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[2] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[1] ;
input \mux_top_inst/algorithm_top_inst/ram_rd_addr[0] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[27] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[26] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[25] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[24] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[23] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[22] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[21] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[20] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[19] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[18] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[17] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[16] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[15] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[14] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[13] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[12] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[11] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[10] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[9] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[8] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[7] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[6] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[5] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[4] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[3] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[2] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[1] ;
input \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[0] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[27] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[26] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[25] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[24] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[23] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[22] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[21] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[20] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[19] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[18] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[17] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[16] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[15] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[14] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[13] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[12] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[11] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[10] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[9] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[8] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[7] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[6] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[5] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[4] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[3] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[2] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[1] ;
input \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[0] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[27] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[26] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[25] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[24] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[23] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[22] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[21] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[20] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[19] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[18] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[17] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[16] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[15] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[14] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[13] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[12] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[11] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[10] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[9] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[8] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[7] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[6] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[5] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[4] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[3] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[2] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[1] ;
input \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[0] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[11] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[10] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[9] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[8] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[7] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[6] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[5] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[4] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[3] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[2] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[1] ;
input \mux_top_inst/algorithm_top_inst/cnt_rx_pix[0] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[27] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[26] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[25] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[24] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[23] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[22] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[21] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[20] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[19] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[18] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[17] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[16] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[15] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[14] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[13] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[12] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[11] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[10] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[9] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[8] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[7] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[6] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[5] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[4] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[3] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[2] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[1] ;
input \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[0] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[255] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[254] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[253] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[252] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[251] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[250] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[249] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[248] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[247] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[246] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[245] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[244] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[243] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[242] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[241] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[240] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[239] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[238] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[237] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[236] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[235] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[234] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[233] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[232] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[231] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[230] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[229] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[228] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[227] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[226] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[225] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[224] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[223] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[222] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[221] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[220] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[219] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[218] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[217] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[216] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[215] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[214] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[213] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[212] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[211] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[210] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[209] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[208] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[207] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[206] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[205] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[204] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[203] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[202] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[201] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[200] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[199] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[198] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[197] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[196] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[195] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[194] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[193] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[192] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[191] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[190] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[189] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[188] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[187] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[186] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[185] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[184] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[183] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[182] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[181] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[180] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[179] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[178] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[177] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[176] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[175] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[174] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[173] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[172] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[171] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[170] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[169] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[168] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[167] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[166] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[165] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[164] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[163] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[162] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[161] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[160] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[159] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[158] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[157] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[156] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[155] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[154] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[153] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[152] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[151] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[150] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[149] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[148] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[147] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[146] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[145] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[144] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[143] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[142] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[141] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[140] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[139] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[138] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[137] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[136] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[135] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[134] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[133] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[132] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[131] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[130] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[129] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[128] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[127] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[126] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[125] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[124] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[123] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[122] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[121] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[120] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[119] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[118] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[117] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[116] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[115] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[114] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[113] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[112] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[111] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[110] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[109] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[108] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[107] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[106] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[105] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[104] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[103] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[102] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[101] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[100] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[99] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[98] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[97] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[96] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[95] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[94] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[93] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[92] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[91] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[90] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[89] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[88] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[87] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[86] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[85] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[84] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[83] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[82] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[81] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[80] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[79] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[78] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[77] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[76] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[75] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[74] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[73] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[72] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[71] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[70] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[69] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[68] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[67] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[66] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[65] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[64] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[63] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[62] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[61] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[60] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[59] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[58] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[57] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[56] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[55] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[54] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[53] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[52] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[51] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[50] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[49] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[48] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[47] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[46] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[45] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[44] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[43] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[42] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[41] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[40] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[39] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[38] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[37] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[36] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[35] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[34] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[33] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[32] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[31] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[30] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[29] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[28] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[27] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[26] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[25] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[24] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[23] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[22] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[21] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[20] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[19] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[18] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[17] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[16] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[15] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[14] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[13] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[12] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[11] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[10] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[9] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[8] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[7] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[6] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[5] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[4] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[3] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[2] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[1] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/dout[0] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[6] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[5] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[4] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[3] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[2] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[1] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ada[0] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[255] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[254] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[253] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[252] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[251] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[250] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[249] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[248] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[247] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[246] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[245] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[244] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[243] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[242] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[241] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[240] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[239] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[238] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[237] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[236] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[235] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[234] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[233] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[232] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[231] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[230] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[229] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[228] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[227] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[226] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[225] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[224] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[223] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[222] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[221] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[220] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[219] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[218] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[217] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[216] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[215] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[214] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[213] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[212] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[211] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[210] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[209] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[208] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[207] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[206] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[205] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[204] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[203] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[202] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[201] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[200] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[199] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[198] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[197] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[196] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[195] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[194] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[193] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[192] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[191] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[190] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[189] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[188] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[187] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[186] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[185] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[184] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[183] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[182] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[181] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[180] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[179] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[178] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[177] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[176] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[175] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[174] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[173] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[172] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[171] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[170] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[169] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[168] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[167] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[166] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[165] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[164] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[163] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[162] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[161] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[160] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[159] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[158] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[157] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[156] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[155] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[154] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[153] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[152] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[151] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[150] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[149] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[148] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[147] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[146] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[145] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[144] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[143] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[142] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[141] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[140] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[139] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[138] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[137] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[136] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[135] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[134] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[133] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[132] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[131] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[130] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[129] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[128] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[127] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[126] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[125] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[124] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[123] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[122] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[121] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[120] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[119] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[118] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[117] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[116] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[115] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[114] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[113] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[112] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[111] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[110] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[109] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[108] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[107] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[106] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[105] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[104] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[103] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[102] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[101] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[100] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[99] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[98] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[97] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[96] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[95] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[94] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[93] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[92] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[91] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[90] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[89] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[88] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[87] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[86] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[85] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[84] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[83] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[82] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[81] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[80] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[79] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[78] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[77] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[76] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[75] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[74] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[73] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[72] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[71] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[70] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[69] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[68] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[67] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[66] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[65] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[64] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[63] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[62] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[61] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[60] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[59] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[58] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[57] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[56] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[55] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[54] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[53] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[52] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[51] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[50] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[49] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[48] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[47] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[46] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[45] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[44] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[43] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[42] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[41] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[40] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[39] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[38] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[37] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[36] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[35] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[34] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[33] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[32] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[31] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[30] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[29] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[28] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[27] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[26] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[25] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[24] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[23] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[22] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[21] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[20] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[19] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[18] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[17] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[16] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[15] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[14] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[13] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[12] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[11] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[10] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[9] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[8] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[7] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[6] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[5] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[4] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[3] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[2] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[1] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/din[0] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[6] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[5] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[4] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[3] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[2] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[1] ;
input \mux_top_inst/algorithm_top_inst/buffer_line/adb[0] ;
input \mux_top_inst/algorithm_top_inst/syn_off0_vs ;
input \mux_top_inst/algorithm_top_inst/coms0_wr_area ;
input \mux_top_inst/algorithm_top_inst/coms1_wr_area ;
input \mux_top_inst/algorithm_top_inst/coms2_wr_area ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.req ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.finish ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.ack ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.data_req ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.req ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.ack ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.dv ;
input \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.finish ;
input \mux_top_inst/algorithm_top_inst/cs_r1 ;
input \mux_top_inst/algorithm_top_inst/cs_r2 ;
input \mux_top_inst/algorithm_top_inst/cs_rise ;
input \mux_top_inst/algorithm_top_inst/ram_rd_en ;
input \mux_top_inst/algorithm_top_inst/ram_wr_en ;
input \mux_top_inst/algorithm_top_inst/buffer_line/clka ;
input \mux_top_inst/algorithm_top_inst/buffer_line/cea ;
input \mux_top_inst/algorithm_top_inst/buffer_line/clkb ;
input \mux_top_inst/algorithm_top_inst/buffer_line/ceb ;
input \mux_top_inst/algorithm_top_inst/buffer_line/oce ;
input \mux_top_inst/algorithm_top_inst/buffer_line/reset ;
input \mux_top_inst/hdmi_rd_inst/ddr_clk ;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[27] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[26] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[25] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[24] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[23] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[22] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[21] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[20] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[19] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[18] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[17] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[16] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[15] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[14] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[13] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[12] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[11] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[10] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[9] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[8] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[7] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/current_buffer_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[28] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[27] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[26] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[25] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[24] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[23] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[22] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[21] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[20] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[19] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[18] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[17] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[16] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[15] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[14] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[13] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[12] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[11] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[10] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[9] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[8] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[7] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[6] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[5] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[4] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[3] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[2] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[1] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[0] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[15] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[14] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[13] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[12] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[11] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[10] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[9] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[8] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[7] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[6] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[5] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[4] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[3] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[2] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[1] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[0] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[255] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[254] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[253] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[252] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[251] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[250] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[249] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[248] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[247] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[246] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[245] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[244] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[243] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[242] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[241] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[240] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[239] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[238] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[237] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[236] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[235] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[234] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[233] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[232] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[231] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[230] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[229] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[228] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[227] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[226] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[225] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[224] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[223] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[222] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[221] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[220] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[219] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[218] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[217] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[216] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[215] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[214] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[213] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[212] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[211] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[210] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[209] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[208] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[207] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[206] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[205] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[204] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[203] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[202] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[201] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[200] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[199] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[198] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[197] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[196] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[195] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[194] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[193] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[192] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[191] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[190] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[189] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[188] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[187] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[186] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[185] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[184] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[183] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[182] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[181] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[180] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[179] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[178] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[177] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[176] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[175] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[174] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[173] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[172] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[171] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[170] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[169] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[168] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[167] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[166] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[165] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[164] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[163] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[162] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[161] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[160] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[159] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[158] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[157] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[156] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[155] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[154] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[153] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[152] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[151] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[150] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[149] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[148] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[147] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[146] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[145] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[144] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[143] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[142] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[141] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[140] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[139] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[138] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[137] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[136] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[135] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[134] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[133] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[132] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[131] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[130] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[129] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[128] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[127] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[126] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[125] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[124] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[123] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[122] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[121] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[120] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[119] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[118] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[117] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[116] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[115] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[114] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[113] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[112] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[111] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[110] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[109] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[108] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[107] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[106] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[105] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[104] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[103] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[102] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[101] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[100] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[99] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[98] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[97] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[96] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[95] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[94] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[93] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[92] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[91] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[90] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[89] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[88] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[87] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[86] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[85] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[84] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[83] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[82] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[81] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[80] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[79] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[78] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[77] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[76] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[75] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[74] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[73] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[72] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[71] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[70] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[69] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[68] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[67] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[66] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[65] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[64] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[63] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[62] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[61] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[60] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[59] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[58] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[57] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[56] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[55] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[54] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[53] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[52] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[51] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[50] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[49] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[48] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[47] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[46] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[45] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[44] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[43] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[42] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[41] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[40] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[39] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[38] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[37] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[36] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[35] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[34] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[33] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[32] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[31] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[30] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[29] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[28] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[27] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[26] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[25] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[24] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[23] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[22] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[21] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[20] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[19] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[18] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[17] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[16] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[15] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[14] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[13] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[12] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[11] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[10] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[9] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[8] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[7] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[6] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[5] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[4] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[3] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[2] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[1] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[0] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[28] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[27] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[26] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[25] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[24] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[23] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[22] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[21] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[20] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[19] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[18] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[17] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[16] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[15] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[14] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[13] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[12] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[11] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[10] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[9] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[8] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[7] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[6] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[5] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[4] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[3] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[2] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[1] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[0] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[15] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[14] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[13] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[12] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[11] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[10] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[9] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[8] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[7] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[6] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[5] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[4] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[3] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[2] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[1] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[0] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[255] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[254] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[253] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[252] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[251] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[250] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[249] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[248] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[247] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[246] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[245] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[244] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[243] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[242] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[241] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[240] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[239] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[238] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[237] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[236] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[235] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[234] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[233] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[232] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[231] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[230] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[229] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[228] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[227] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[226] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[225] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[224] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[223] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[222] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[221] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[220] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[219] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[218] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[217] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[216] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[215] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[214] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[213] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[212] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[211] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[210] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[209] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[208] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[207] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[206] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[205] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[204] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[203] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[202] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[201] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[200] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[199] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[198] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[197] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[196] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[195] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[194] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[193] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[192] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[191] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[190] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[189] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[188] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[187] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[186] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[185] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[184] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[183] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[182] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[181] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[180] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[179] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[178] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[177] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[176] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[175] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[174] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[173] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[172] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[171] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[170] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[169] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[168] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[167] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[166] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[165] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[164] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[163] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[162] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[161] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[160] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[159] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[158] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[157] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[156] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[155] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[154] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[153] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[152] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[151] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[150] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[149] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[148] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[147] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[146] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[145] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[144] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[143] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[142] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[141] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[140] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[139] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[138] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[137] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[136] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[135] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[134] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[133] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[132] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[131] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[130] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[129] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[128] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[127] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[126] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[125] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[124] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[123] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[122] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[121] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[120] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[119] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[118] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[117] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[116] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[115] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[114] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[113] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[112] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[111] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[110] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[109] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[108] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[107] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[106] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[105] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[104] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[103] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[102] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[101] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[100] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[99] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[98] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[97] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[96] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[95] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[94] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[93] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[92] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[91] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[90] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[89] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[88] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[87] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[86] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[85] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[84] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[83] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[82] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[81] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[80] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[79] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[78] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[77] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[76] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[75] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[74] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[73] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[72] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[71] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[70] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[69] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[68] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[67] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[66] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[65] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[64] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[63] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[62] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[61] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[60] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[59] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[58] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[57] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[56] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[55] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[54] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[53] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[52] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[51] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[50] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[49] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[48] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[47] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[46] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[45] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[44] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[43] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[42] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[41] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[40] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[39] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[38] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[37] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[36] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[35] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[34] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[33] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[32] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[31] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[30] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[29] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[28] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[27] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[26] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[25] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[24] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[23] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[22] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[21] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[20] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[19] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[18] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[17] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[16] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[15] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[14] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[13] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[12] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[11] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[10] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[9] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[8] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[7] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[6] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[5] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[4] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[3] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[2] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[1] ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[0] ;
wire \mux_top_inst/algorithm_top_inst/time_out[19] ;
wire \mux_top_inst/algorithm_top_inst/time_out[18] ;
wire \mux_top_inst/algorithm_top_inst/time_out[17] ;
wire \mux_top_inst/algorithm_top_inst/time_out[16] ;
wire \mux_top_inst/algorithm_top_inst/time_out[15] ;
wire \mux_top_inst/algorithm_top_inst/time_out[14] ;
wire \mux_top_inst/algorithm_top_inst/time_out[13] ;
wire \mux_top_inst/algorithm_top_inst/time_out[12] ;
wire \mux_top_inst/algorithm_top_inst/time_out[11] ;
wire \mux_top_inst/algorithm_top_inst/time_out[10] ;
wire \mux_top_inst/algorithm_top_inst/time_out[9] ;
wire \mux_top_inst/algorithm_top_inst/time_out[8] ;
wire \mux_top_inst/algorithm_top_inst/time_out[7] ;
wire \mux_top_inst/algorithm_top_inst/time_out[6] ;
wire \mux_top_inst/algorithm_top_inst/time_out[5] ;
wire \mux_top_inst/algorithm_top_inst/time_out[4] ;
wire \mux_top_inst/algorithm_top_inst/time_out[3] ;
wire \mux_top_inst/algorithm_top_inst/time_out[2] ;
wire \mux_top_inst/algorithm_top_inst/time_out[1] ;
wire \mux_top_inst/algorithm_top_inst/time_out[0] ;
wire \mux_top_inst/algorithm_top_inst/cs[7] ;
wire \mux_top_inst/algorithm_top_inst/cs[6] ;
wire \mux_top_inst/algorithm_top_inst/cs[5] ;
wire \mux_top_inst/algorithm_top_inst/cs[4] ;
wire \mux_top_inst/algorithm_top_inst/cs[3] ;
wire \mux_top_inst/algorithm_top_inst/cs[2] ;
wire \mux_top_inst/algorithm_top_inst/cs[1] ;
wire \mux_top_inst/algorithm_top_inst/cs[0] ;
wire \mux_top_inst/algorithm_top_inst/cmos_cnt[4] ;
wire \mux_top_inst/algorithm_top_inst/cmos_cnt[3] ;
wire \mux_top_inst/algorithm_top_inst/cmos_cnt[2] ;
wire \mux_top_inst/algorithm_top_inst/cmos_cnt[1] ;
wire \mux_top_inst/algorithm_top_inst/cmos_cnt[0] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[10] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[9] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[8] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[7] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[6] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[5] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[4] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[3] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[2] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[1] ;
wire \mux_top_inst/algorithm_top_inst/line_cnt[0] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[255] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[254] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[253] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[252] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[251] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[250] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[249] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[248] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[247] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[246] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[245] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[244] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[243] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[242] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[241] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[240] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[239] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[238] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[237] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[236] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[235] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[234] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[233] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[232] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[231] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[230] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[229] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[228] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[227] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[226] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[225] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[224] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[223] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[222] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[221] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[220] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[219] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[218] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[217] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[216] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[215] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[214] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[213] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[212] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[211] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[210] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[209] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[208] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[207] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[206] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[205] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[204] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[203] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[202] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[201] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[200] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[199] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[198] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[197] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[196] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[195] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[194] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[193] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[192] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[191] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[190] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[189] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[188] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[187] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[186] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[185] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[184] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[183] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[182] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[181] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[180] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[179] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[178] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[177] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[176] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[175] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[174] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[173] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[172] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[171] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[170] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[169] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[168] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[167] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[166] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[165] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[164] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[163] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[162] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[161] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[160] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[159] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[158] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[157] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[156] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[155] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[154] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[153] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[152] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[151] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[150] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[149] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[148] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[147] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[146] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[145] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[144] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[143] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[142] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[141] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[140] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[139] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[138] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[137] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[136] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[135] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[134] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[133] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[132] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[131] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[130] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[129] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[128] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[127] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[126] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[125] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[124] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[123] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[122] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[121] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[120] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[119] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[118] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[117] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[116] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[115] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[114] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[113] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[112] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[111] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[110] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[109] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[108] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[107] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[106] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[105] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[104] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[103] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[102] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[101] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[100] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[99] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[98] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[97] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[96] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[95] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[94] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[93] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[92] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[91] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[90] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[89] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[88] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[87] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[86] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[85] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[84] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[83] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[82] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[81] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[80] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[79] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[78] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[77] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[76] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[75] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[74] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[73] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[72] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[71] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[70] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[69] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[68] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[67] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[66] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[65] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[64] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[63] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[62] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[61] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[60] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[59] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[58] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[57] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[56] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[55] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[54] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[53] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[52] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[51] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[50] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[49] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[48] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[47] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[46] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[45] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[44] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[43] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[42] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[41] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[40] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[39] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[38] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[37] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[36] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[35] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[34] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[33] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[32] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[31] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[30] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[29] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[28] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[27] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[26] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[25] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[24] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[23] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[22] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[21] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[20] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[19] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[18] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[17] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[16] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[15] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[14] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[13] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[12] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[11] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[10] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[9] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[8] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[7] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[6] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[5] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[4] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[3] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[2] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[1] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_data[0] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[255] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[254] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[253] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[252] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[251] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[250] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[249] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[248] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[247] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[246] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[245] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[244] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[243] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[242] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[241] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[240] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[239] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[238] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[237] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[236] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[235] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[234] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[233] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[232] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[231] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[230] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[229] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[228] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[227] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[226] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[225] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[224] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[223] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[222] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[221] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[220] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[219] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[218] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[217] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[216] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[215] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[214] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[213] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[212] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[211] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[210] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[209] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[208] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[207] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[206] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[205] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[204] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[203] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[202] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[201] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[200] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[199] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[198] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[197] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[196] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[195] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[194] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[193] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[192] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[191] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[190] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[189] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[188] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[187] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[186] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[185] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[184] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[183] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[182] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[181] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[180] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[179] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[178] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[177] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[176] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[175] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[174] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[173] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[172] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[171] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[170] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[169] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[168] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[167] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[166] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[165] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[164] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[163] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[162] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[161] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[160] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[159] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[158] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[157] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[156] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[155] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[154] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[153] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[152] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[151] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[150] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[149] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[148] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[147] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[146] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[145] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[144] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[143] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[142] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[141] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[140] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[139] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[138] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[137] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[136] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[135] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[134] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[133] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[132] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[131] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[130] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[129] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[128] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[127] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[126] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[125] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[124] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[123] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[122] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[121] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[120] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[119] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[118] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[117] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[116] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[115] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[114] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[113] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[112] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[111] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[110] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[109] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[108] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[107] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[106] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[105] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[104] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[103] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[102] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[101] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[100] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[99] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[98] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[97] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[96] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[95] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[94] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[93] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[92] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[91] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[90] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[89] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[88] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[87] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[86] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[85] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[84] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[83] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[82] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[81] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[80] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[79] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[78] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[77] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[76] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[75] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[74] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[73] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[72] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[71] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[70] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[69] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[68] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[67] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[66] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[65] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[64] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[63] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[62] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[61] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[60] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[59] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[58] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[57] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[56] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[55] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[54] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[53] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[52] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[51] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[50] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[49] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[48] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[47] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[46] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[45] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[44] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[43] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[42] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[41] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[40] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[39] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[38] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[37] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[36] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[35] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[34] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[33] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[32] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[31] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[30] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[29] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[28] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[27] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[26] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[25] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[24] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[23] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[22] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[21] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[20] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[19] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[18] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[17] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[16] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[15] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[14] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[13] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[12] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[11] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[10] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[9] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[8] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[7] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[6] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[5] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[4] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[3] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[2] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[1] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_data[0] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[27] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[26] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[25] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[24] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[23] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[22] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[21] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[20] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[19] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[18] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[17] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[16] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[15] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[14] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[13] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[12] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[11] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[10] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[9] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[8] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[7] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/cmos0_rd_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[27] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[26] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[25] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[24] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[23] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[22] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[21] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[20] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[19] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[18] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[17] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[16] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[15] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[14] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[13] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[12] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[11] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[10] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[9] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[8] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[7] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/cmos1_rd_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[27] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[26] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[25] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[24] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[23] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[22] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[21] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[20] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[19] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[18] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[17] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[16] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[15] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[14] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[13] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[12] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[11] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[10] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[9] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[8] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[7] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/cmos2_rd_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[11] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[10] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[9] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[8] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[7] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[6] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[5] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[4] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[3] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[2] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[1] ;
wire \mux_top_inst/algorithm_top_inst/cnt_rx_pix[0] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[27] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[26] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[25] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[24] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[23] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[22] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[21] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[20] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[19] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[18] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[17] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[16] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[15] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[14] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[13] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[12] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[11] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[10] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[9] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[8] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[7] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[6] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[5] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[4] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[3] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[2] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[1] ;
wire \mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[0] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[255] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[254] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[253] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[252] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[251] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[250] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[249] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[248] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[247] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[246] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[245] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[244] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[243] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[242] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[241] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[240] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[239] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[238] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[237] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[236] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[235] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[234] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[233] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[232] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[231] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[230] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[229] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[228] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[227] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[226] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[225] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[224] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[223] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[222] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[221] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[220] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[219] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[218] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[217] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[216] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[215] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[214] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[213] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[212] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[211] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[210] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[209] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[208] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[207] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[206] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[205] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[204] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[203] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[202] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[201] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[200] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[199] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[198] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[197] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[196] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[195] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[194] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[193] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[192] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[191] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[190] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[189] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[188] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[187] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[186] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[185] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[184] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[183] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[182] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[181] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[180] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[179] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[178] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[177] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[176] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[175] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[174] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[173] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[172] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[171] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[170] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[169] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[168] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[167] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[166] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[165] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[164] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[163] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[162] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[161] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[160] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[159] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[158] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[157] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[156] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[155] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[154] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[153] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[152] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[151] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[150] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[149] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[148] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[147] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[146] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[145] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[144] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[143] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[142] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[141] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[140] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[139] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[138] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[137] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[136] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[135] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[134] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[133] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[132] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[131] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[130] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[129] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[128] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[127] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[126] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[125] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[124] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[123] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[122] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[121] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[120] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[119] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[118] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[117] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[116] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[115] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[114] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[113] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[112] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[111] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[110] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[109] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[108] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[107] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[106] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[105] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[104] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[103] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[102] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[101] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[100] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[99] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[98] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[97] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[96] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[95] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[94] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[93] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[92] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[91] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[90] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[89] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[88] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[87] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[86] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[85] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[84] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[83] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[82] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[81] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[80] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[79] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[78] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[77] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[76] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[75] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[74] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[73] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[72] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[71] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[70] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[69] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[68] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[67] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[66] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[65] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[64] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[63] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[62] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[61] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[60] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[59] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[58] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[57] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[56] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[55] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[54] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[53] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[52] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[51] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[50] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[49] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[48] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[47] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[46] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[45] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[44] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[43] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[42] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[41] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[40] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[39] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[38] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[37] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[36] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[35] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[34] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[33] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[32] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[31] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[30] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[29] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[28] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[27] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[26] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[25] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[24] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[23] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[22] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[21] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[20] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[19] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[18] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[17] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[16] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[15] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[14] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[13] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[12] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[11] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[10] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[9] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[8] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[7] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[6] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[5] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[4] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[3] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[2] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[1] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/dout[0] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[6] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[5] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[4] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[3] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[2] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[1] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ada[0] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[255] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[254] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[253] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[252] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[251] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[250] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[249] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[248] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[247] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[246] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[245] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[244] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[243] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[242] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[241] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[240] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[239] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[238] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[237] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[236] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[235] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[234] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[233] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[232] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[231] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[230] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[229] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[228] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[227] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[226] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[225] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[224] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[223] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[222] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[221] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[220] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[219] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[218] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[217] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[216] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[215] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[214] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[213] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[212] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[211] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[210] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[209] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[208] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[207] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[206] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[205] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[204] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[203] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[202] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[201] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[200] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[199] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[198] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[197] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[196] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[195] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[194] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[193] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[192] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[191] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[190] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[189] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[188] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[187] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[186] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[185] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[184] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[183] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[182] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[181] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[180] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[179] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[178] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[177] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[176] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[175] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[174] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[173] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[172] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[171] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[170] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[169] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[168] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[167] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[166] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[165] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[164] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[163] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[162] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[161] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[160] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[159] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[158] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[157] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[156] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[155] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[154] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[153] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[152] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[151] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[150] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[149] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[148] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[147] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[146] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[145] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[144] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[143] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[142] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[141] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[140] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[139] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[138] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[137] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[136] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[135] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[134] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[133] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[132] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[131] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[130] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[129] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[128] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[127] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[126] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[125] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[124] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[123] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[122] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[121] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[120] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[119] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[118] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[117] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[116] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[115] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[114] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[113] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[112] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[111] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[110] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[109] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[108] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[107] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[106] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[105] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[104] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[103] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[102] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[101] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[100] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[99] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[98] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[97] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[96] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[95] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[94] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[93] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[92] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[91] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[90] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[89] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[88] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[87] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[86] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[85] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[84] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[83] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[82] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[81] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[80] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[79] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[78] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[77] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[76] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[75] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[74] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[73] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[72] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[71] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[70] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[69] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[68] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[67] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[66] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[65] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[64] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[63] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[62] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[61] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[60] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[59] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[58] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[57] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[56] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[55] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[54] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[53] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[52] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[51] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[50] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[49] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[48] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[47] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[46] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[45] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[44] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[43] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[42] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[41] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[40] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[39] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[38] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[37] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[36] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[35] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[34] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[33] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[32] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[31] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[30] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[29] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[28] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[27] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[26] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[25] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[24] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[23] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[22] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[21] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[20] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[19] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[18] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[17] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[16] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[15] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[14] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[13] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[12] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[11] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[10] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[9] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[8] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[7] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[6] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[5] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[4] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[3] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[2] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[1] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/din[0] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[6] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[5] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[4] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[3] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[2] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[1] ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/adb[0] ;
wire \mux_top_inst/algorithm_top_inst/syn_off0_vs ;
wire \mux_top_inst/algorithm_top_inst/coms0_wr_area ;
wire \mux_top_inst/algorithm_top_inst/coms1_wr_area ;
wire \mux_top_inst/algorithm_top_inst/coms2_wr_area ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.req ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.finish ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.ack ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.data_req ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.req ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.ack ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.dv ;
wire \mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.finish ;
wire \mux_top_inst/algorithm_top_inst/cs_r1 ;
wire \mux_top_inst/algorithm_top_inst/cs_r2 ;
wire \mux_top_inst/algorithm_top_inst/cs_rise ;
wire \mux_top_inst/algorithm_top_inst/ram_rd_en ;
wire \mux_top_inst/algorithm_top_inst/ram_wr_en ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/clka ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/cea ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/clkb ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/ceb ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/oce ;
wire \mux_top_inst/algorithm_top_inst/buffer_line/reset ;
wire \mux_top_inst/hdmi_rd_inst/ddr_clk ;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\mux_top_inst/algorithm_top_inst/cs[7] ,\mux_top_inst/algorithm_top_inst/cs[6] ,\mux_top_inst/algorithm_top_inst/cs[5] ,\mux_top_inst/algorithm_top_inst/cs[4] ,\mux_top_inst/algorithm_top_inst/cs[3] ,\mux_top_inst/algorithm_top_inst/cs[2] ,\mux_top_inst/algorithm_top_inst/cs[1] ,\mux_top_inst/algorithm_top_inst/cs[0] ,\mux_top_inst/algorithm_top_inst/line_cnt[10] ,\mux_top_inst/algorithm_top_inst/line_cnt[9] ,\mux_top_inst/algorithm_top_inst/line_cnt[8] ,\mux_top_inst/algorithm_top_inst/line_cnt[7] ,\mux_top_inst/algorithm_top_inst/line_cnt[6] ,\mux_top_inst/algorithm_top_inst/line_cnt[5] ,\mux_top_inst/algorithm_top_inst/line_cnt[4] ,\mux_top_inst/algorithm_top_inst/line_cnt[3] ,\mux_top_inst/algorithm_top_inst/line_cnt[2] ,\mux_top_inst/algorithm_top_inst/line_cnt[1] ,\mux_top_inst/algorithm_top_inst/line_cnt[0] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[11] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[10] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[9] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[8] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[7] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[6] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[5] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[4] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[3] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[2] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[1] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[0] ,\mux_top_inst/algorithm_top_inst/cs_rise ,\mux_top_inst/algorithm_top_inst/ram_wr_en ,\mux_top_inst/algorithm_top_inst/ram_rd_en }),
    .data_i({\mux_top_inst/algorithm_top_inst/current_buffer_addr[27] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[26] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[25] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[24] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[23] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[22] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[21] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[20] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[19] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[18] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[17] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[16] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[15] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[14] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[13] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[12] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[11] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[10] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[9] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[8] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[7] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[6] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[5] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[4] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[3] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[2] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[1] ,\mux_top_inst/algorithm_top_inst/current_buffer_addr[0] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[28] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[27] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[26] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[25] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[24] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[23] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[22] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[21] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[20] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[19] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[18] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[17] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[16] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[15] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[14] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[13] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[12] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[11] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[10] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[9] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[8] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[7] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[6] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[5] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[4] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[3] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[2] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[1] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.addr[0] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[15] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[14] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[13] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[12] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[11] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[10] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[9] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[8] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[7] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[6] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[5] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[4] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[3] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[2] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[1] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.len[0] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[255] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[254] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[253] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[252] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[251] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[250] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[249] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[248] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[247] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[246] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[245] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[244] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[243] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[242] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[241] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[240] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[239] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[238] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[237] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[236] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[235] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[234] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[233] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[232] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[231] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[230] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[229] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[228] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[227] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[226] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[225] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[224] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[223] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[222] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[221] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[220] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[219] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[218] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[217] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[216] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[215] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[214] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[213] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[212] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[211] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[210] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[209] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[208] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[207] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[206] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[205] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[204] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[203] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[202] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[201] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[200] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[199] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[198] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[197] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[196] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[195] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[194] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[193] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[192] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[191] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[190] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[189] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[188] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[187] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[186] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[185] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[184] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[183] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[182] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[181] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[180] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[179] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[178] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[177] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[176] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[175] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[174] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[173] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[172] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[171] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[170] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[169] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[168] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[167] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[166] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[165] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[164] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[163] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[162] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[161] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[160] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[159] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[158] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[157] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[156] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[155] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[154] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[153] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[152] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[151] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[150] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[149] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[148] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[147] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[146] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[145] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[144] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[143] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[142] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[141] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[140] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[139] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[138] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[137] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[136] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[135] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[134] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[133] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[132] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[131] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[130] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[129] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[128] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[127] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[126] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[125] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[124] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[123] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[122] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[121] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[120] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[119] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[118] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[117] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[116] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[115] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[114] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[113] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[112] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[111] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[110] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[109] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[108] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[107] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[106] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[105] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[104] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[103] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[102] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[101] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[100] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[99] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[98] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[97] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[96] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[95] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[94] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[93] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[92] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[91] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[90] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[89] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[88] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[87] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[86] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[85] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[84] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[83] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[82] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[81] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[80] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[79] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[78] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[77] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[76] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[75] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[74] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[73] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[72] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[71] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[70] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[69] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[68] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[67] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[66] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[65] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[64] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[63] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[62] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[61] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[60] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[59] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[58] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[57] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[56] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[55] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[54] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[53] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[52] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[51] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[50] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[49] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[48] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[47] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[46] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[45] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[44] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[43] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[42] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[41] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[40] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[39] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[38] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[37] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[36] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[35] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[34] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[33] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[32] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[31] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[30] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[29] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[28] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[27] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[26] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[25] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[24] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[23] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[22] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[21] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[20] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[19] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[18] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[17] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[16] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[15] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[14] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[13] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[12] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[11] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[10] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[9] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[8] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[7] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[6] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[5] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[4] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[3] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[2] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[1] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.data[0] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[28] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[27] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[26] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[25] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[24] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[23] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[22] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[21] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[20] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[19] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[18] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[17] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[16] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[15] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[14] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[13] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[12] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[11] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[10] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[9] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[8] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[7] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[6] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[5] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[4] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[3] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[2] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[1] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.addr[0] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[15] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[14] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[13] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[12] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[11] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[10] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[9] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[8] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[7] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[6] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[5] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[4] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[3] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[2] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[1] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.len[0] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[255] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[254] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[253] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[252] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[251] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[250] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[249] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[248] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[247] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[246] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[245] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[244] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[243] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[242] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[241] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[240] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[239] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[238] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[237] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[236] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[235] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[234] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[233] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[232] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[231] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[230] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[229] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[228] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[227] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[226] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[225] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[224] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[223] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[222] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[221] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[220] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[219] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[218] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[217] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[216] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[215] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[214] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[213] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[212] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[211] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[210] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[209] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[208] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[207] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[206] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[205] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[204] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[203] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[202] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[201] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[200] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[199] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[198] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[197] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[196] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[195] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[194] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[193] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[192] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[191] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[190] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[189] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[188] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[187] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[186] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[185] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[184] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[183] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[182] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[181] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[180] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[179] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[178] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[177] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[176] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[175] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[174] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[173] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[172] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[171] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[170] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[169] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[168] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[167] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[166] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[165] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[164] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[163] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[162] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[161] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[160] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[159] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[158] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[157] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[156] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[155] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[154] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[153] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[152] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[151] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[150] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[149] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[148] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[147] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[146] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[145] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[144] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[143] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[142] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[141] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[140] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[139] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[138] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[137] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[136] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[135] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[134] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[133] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[132] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[131] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[130] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[129] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[128] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[127] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[126] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[125] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[124] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[123] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[122] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[121] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[120] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[119] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[118] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[117] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[116] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[115] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[114] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[113] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[112] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[111] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[110] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[109] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[108] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[107] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[106] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[105] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[104] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[103] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[102] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[101] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[100] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[99] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[98] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[97] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[96] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[95] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[94] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[93] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[92] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[91] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[90] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[89] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[88] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[87] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[86] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[85] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[84] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[83] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[82] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[81] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[80] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[79] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[78] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[77] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[76] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[75] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[74] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[73] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[72] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[71] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[70] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[69] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[68] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[67] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[66] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[65] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[64] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[63] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[62] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[61] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[60] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[59] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[58] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[57] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[56] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[55] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[54] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[53] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[52] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[51] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[50] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[49] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[48] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[47] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[46] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[45] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[44] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[43] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[42] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[41] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[40] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[39] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[38] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[37] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[36] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[35] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[34] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[33] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[32] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[31] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[30] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[29] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[28] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[27] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[26] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[25] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[24] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[23] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[22] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[21] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[20] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[19] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[18] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[17] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[16] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[15] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[14] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[13] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[12] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[11] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[10] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[9] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[8] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[7] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[6] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[5] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[4] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[3] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[2] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[1] ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.data[0] ,\mux_top_inst/algorithm_top_inst/time_out[19] ,\mux_top_inst/algorithm_top_inst/time_out[18] ,\mux_top_inst/algorithm_top_inst/time_out[17] ,\mux_top_inst/algorithm_top_inst/time_out[16] ,\mux_top_inst/algorithm_top_inst/time_out[15] ,\mux_top_inst/algorithm_top_inst/time_out[14] ,\mux_top_inst/algorithm_top_inst/time_out[13] ,\mux_top_inst/algorithm_top_inst/time_out[12] ,\mux_top_inst/algorithm_top_inst/time_out[11] ,\mux_top_inst/algorithm_top_inst/time_out[10] ,\mux_top_inst/algorithm_top_inst/time_out[9] ,\mux_top_inst/algorithm_top_inst/time_out[8] ,\mux_top_inst/algorithm_top_inst/time_out[7] ,\mux_top_inst/algorithm_top_inst/time_out[6] ,\mux_top_inst/algorithm_top_inst/time_out[5] ,\mux_top_inst/algorithm_top_inst/time_out[4] ,\mux_top_inst/algorithm_top_inst/time_out[3] ,\mux_top_inst/algorithm_top_inst/time_out[2] ,\mux_top_inst/algorithm_top_inst/time_out[1] ,\mux_top_inst/algorithm_top_inst/time_out[0] ,\mux_top_inst/algorithm_top_inst/cs[7] ,\mux_top_inst/algorithm_top_inst/cs[6] ,\mux_top_inst/algorithm_top_inst/cs[5] ,\mux_top_inst/algorithm_top_inst/cs[4] ,\mux_top_inst/algorithm_top_inst/cs[3] ,\mux_top_inst/algorithm_top_inst/cs[2] ,\mux_top_inst/algorithm_top_inst/cs[1] ,\mux_top_inst/algorithm_top_inst/cs[0] ,\mux_top_inst/algorithm_top_inst/cmos_cnt[4] ,\mux_top_inst/algorithm_top_inst/cmos_cnt[3] ,\mux_top_inst/algorithm_top_inst/cmos_cnt[2] ,\mux_top_inst/algorithm_top_inst/cmos_cnt[1] ,\mux_top_inst/algorithm_top_inst/cmos_cnt[0] ,\mux_top_inst/algorithm_top_inst/line_cnt[10] ,\mux_top_inst/algorithm_top_inst/line_cnt[9] ,\mux_top_inst/algorithm_top_inst/line_cnt[8] ,\mux_top_inst/algorithm_top_inst/line_cnt[7] ,\mux_top_inst/algorithm_top_inst/line_cnt[6] ,\mux_top_inst/algorithm_top_inst/line_cnt[5] ,\mux_top_inst/algorithm_top_inst/line_cnt[4] ,\mux_top_inst/algorithm_top_inst/line_cnt[3] ,\mux_top_inst/algorithm_top_inst/line_cnt[2] ,\mux_top_inst/algorithm_top_inst/line_cnt[1] ,\mux_top_inst/algorithm_top_inst/line_cnt[0] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[255] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[254] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[253] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[252] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[251] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[250] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[249] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[248] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[247] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[246] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[245] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[244] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[243] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[242] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[241] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[240] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[239] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[238] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[237] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[236] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[235] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[234] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[233] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[232] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[231] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[230] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[229] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[228] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[227] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[226] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[225] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[224] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[223] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[222] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[221] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[220] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[219] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[218] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[217] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[216] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[215] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[214] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[213] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[212] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[211] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[210] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[209] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[208] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[207] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[206] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[205] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[204] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[203] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[202] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[201] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[200] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[199] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[198] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[197] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[196] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[195] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[194] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[193] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[192] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[191] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[190] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[189] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[188] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[187] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[186] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[185] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[184] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[183] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[182] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[181] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[180] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[179] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[178] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[177] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[176] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[175] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[174] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[173] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[172] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[171] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[170] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[169] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[168] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[167] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[166] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[165] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[164] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[163] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[162] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[161] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[160] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[159] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[158] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[157] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[156] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[155] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[154] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[153] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[152] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[151] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[150] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[149] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[148] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[147] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[146] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[145] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[144] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[143] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[142] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[141] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[140] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[139] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[138] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[137] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[136] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[135] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[134] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[133] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[132] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[131] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[130] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[129] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[128] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[127] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[126] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[125] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[124] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[123] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[122] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[121] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[120] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[119] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[118] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[117] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[116] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[115] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[114] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[113] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[112] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[111] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[110] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[109] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[108] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[107] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[106] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[105] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[104] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[103] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[102] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[101] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[100] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[99] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[98] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[97] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[96] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[95] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[94] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[93] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[92] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[91] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[90] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[89] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[88] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[87] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[86] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[85] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[84] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[83] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[82] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[81] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[80] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[79] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[78] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[77] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[76] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[75] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[74] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[73] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[72] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[71] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[70] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[69] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[68] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[67] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[66] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[65] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[64] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[63] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[62] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[61] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[60] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[59] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[58] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[57] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[56] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[55] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[54] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[53] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[52] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[51] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[50] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[49] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[48] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[47] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[46] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[45] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[44] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[43] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[42] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[41] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[40] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[39] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[38] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[37] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[36] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[35] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[34] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[33] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[32] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[31] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[30] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[29] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[28] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[27] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[26] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[25] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[24] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[23] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[22] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[21] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[20] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[19] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[18] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[17] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[16] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[15] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[14] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[13] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[12] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[11] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[10] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[9] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[8] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[7] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[6] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[5] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[4] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[3] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[2] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[1] ,\mux_top_inst/algorithm_top_inst/ram_rd_data[0] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[255] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[254] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[253] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[252] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[251] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[250] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[249] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[248] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[247] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[246] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[245] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[244] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[243] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[242] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[241] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[240] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[239] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[238] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[237] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[236] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[235] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[234] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[233] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[232] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[231] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[230] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[229] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[228] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[227] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[226] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[225] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[224] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[223] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[222] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[221] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[220] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[219] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[218] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[217] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[216] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[215] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[214] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[213] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[212] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[211] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[210] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[209] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[208] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[207] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[206] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[205] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[204] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[203] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[202] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[201] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[200] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[199] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[198] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[197] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[196] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[195] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[194] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[193] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[192] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[191] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[190] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[189] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[188] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[187] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[186] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[185] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[184] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[183] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[182] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[181] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[180] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[179] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[178] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[177] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[176] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[175] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[174] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[173] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[172] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[171] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[170] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[169] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[168] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[167] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[166] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[165] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[164] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[163] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[162] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[161] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[160] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[159] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[158] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[157] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[156] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[155] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[154] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[153] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[152] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[151] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[150] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[149] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[148] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[147] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[146] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[145] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[144] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[143] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[142] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[141] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[140] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[139] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[138] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[137] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[136] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[135] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[134] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[133] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[132] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[131] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[130] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[129] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[128] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[127] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[126] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[125] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[124] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[123] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[122] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[121] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[120] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[119] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[118] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[117] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[116] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[115] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[114] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[113] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[112] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[111] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[110] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[109] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[108] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[107] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[106] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[105] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[104] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[103] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[102] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[101] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[100] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[99] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[98] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[97] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[96] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[95] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[94] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[93] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[92] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[91] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[90] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[89] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[88] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[87] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[86] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[85] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[84] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[83] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[82] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[81] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[80] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[79] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[78] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[77] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[76] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[75] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[74] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[73] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[72] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[71] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[70] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[69] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[68] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[67] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[66] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[65] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[64] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[63] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[62] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[61] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[60] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[59] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[58] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[57] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[56] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[55] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[54] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[53] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[52] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[51] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[50] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[49] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[48] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[47] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[46] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[45] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[44] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[43] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[42] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[41] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[40] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[39] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[38] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[37] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[36] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[35] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[34] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[33] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[32] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[31] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[30] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[29] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[28] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[27] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[26] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[25] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[24] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[23] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[22] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[21] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[20] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[19] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[18] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[17] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[16] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[15] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[14] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[13] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[12] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[11] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[10] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[9] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[8] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[7] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[6] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[5] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[4] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[3] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[2] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[1] ,\mux_top_inst/algorithm_top_inst/ram_wr_data[0] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[6] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[5] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[4] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[3] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[2] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[1] ,\mux_top_inst/algorithm_top_inst/ram_wr_addr[0] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[6] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[5] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[4] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[3] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[2] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[1] ,\mux_top_inst/algorithm_top_inst/ram_rd_addr[0] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[27] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[26] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[25] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[24] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[23] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[22] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[21] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[20] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[19] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[18] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[17] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[16] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[15] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[14] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[13] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[12] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[11] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[10] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[9] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[8] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[7] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[6] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[5] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[4] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[3] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[2] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[1] ,\mux_top_inst/algorithm_top_inst/cmos0_rd_addr[0] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[27] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[26] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[25] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[24] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[23] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[22] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[21] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[20] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[19] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[18] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[17] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[16] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[15] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[14] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[13] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[12] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[11] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[10] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[9] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[8] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[7] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[6] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[5] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[4] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[3] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[2] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[1] ,\mux_top_inst/algorithm_top_inst/cmos1_rd_addr[0] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[27] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[26] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[25] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[24] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[23] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[22] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[21] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[20] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[19] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[18] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[17] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[16] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[15] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[14] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[13] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[12] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[11] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[10] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[9] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[8] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[7] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[6] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[5] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[4] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[3] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[2] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[1] ,\mux_top_inst/algorithm_top_inst/cmos2_rd_addr[0] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[11] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[10] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[9] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[8] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[7] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[6] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[5] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[4] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[3] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[2] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[1] ,\mux_top_inst/algorithm_top_inst/cnt_rx_pix[0] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[27] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[26] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[25] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[24] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[23] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[22] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[21] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[20] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[19] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[18] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[17] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[16] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[15] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[14] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[13] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[12] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[11] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[10] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[9] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[8] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[7] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[6] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[5] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[4] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[3] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[2] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[1] ,\mux_top_inst/algorithm_top_inst/ddr_wr_init_addr[0] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[255] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[254] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[253] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[252] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[251] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[250] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[249] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[248] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[247] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[246] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[245] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[244] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[243] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[242] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[241] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[240] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[239] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[238] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[237] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[236] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[235] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[234] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[233] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[232] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[231] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[230] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[229] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[228] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[227] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[226] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[225] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[224] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[223] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[222] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[221] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[220] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[219] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[218] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[217] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[216] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[215] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[214] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[213] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[212] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[211] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[210] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[209] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[208] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[207] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[206] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[205] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[204] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[203] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[202] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[201] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[200] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[199] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[198] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[197] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[196] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[195] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[194] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[193] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[192] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[191] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[190] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[189] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[188] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[187] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[186] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[185] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[184] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[183] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[182] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[181] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[180] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[179] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[178] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[177] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[176] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[175] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[174] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[173] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[172] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[171] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[170] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[169] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[168] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[167] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[166] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[165] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[164] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[163] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[162] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[161] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[160] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[159] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[158] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[157] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[156] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[155] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[154] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[153] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[152] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[151] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[150] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[149] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[148] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[147] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[146] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[145] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[144] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[143] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[142] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[141] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[140] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[139] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[138] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[137] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[136] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[135] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[134] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[133] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[132] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[131] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[130] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[129] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[128] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[127] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[126] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[125] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[124] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[123] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[122] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[121] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[120] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[119] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[118] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[117] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[116] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[115] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[114] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[113] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[112] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[111] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[110] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[109] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[108] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[107] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[106] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[105] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[104] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[103] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[102] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[101] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[100] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[99] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[98] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[97] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[96] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[95] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[94] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[93] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[92] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[91] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[90] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[89] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[88] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[87] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[86] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[85] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[84] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[83] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[82] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[81] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[80] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[79] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[78] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[77] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[76] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[75] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[74] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[73] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[72] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[71] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[70] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[69] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[68] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[67] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[66] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[65] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[64] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[63] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[62] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[61] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[60] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[59] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[58] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[57] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[56] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[55] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[54] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[53] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[52] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[51] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[50] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[49] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[48] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[47] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[46] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[45] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[44] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[43] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[42] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[41] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[40] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[39] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[38] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[37] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[36] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[35] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[34] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[33] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[32] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[31] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[30] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[29] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[28] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[27] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[26] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[25] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[24] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[23] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[22] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[21] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[20] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[19] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[18] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[17] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[16] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[15] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[14] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[13] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[12] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[11] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[10] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[9] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[8] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[7] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[6] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[5] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[4] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[3] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[2] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[1] ,\mux_top_inst/algorithm_top_inst/buffer_line/dout[0] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[6] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[5] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[4] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[3] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[2] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[1] ,\mux_top_inst/algorithm_top_inst/buffer_line/ada[0] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[255] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[254] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[253] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[252] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[251] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[250] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[249] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[248] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[247] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[246] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[245] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[244] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[243] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[242] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[241] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[240] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[239] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[238] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[237] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[236] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[235] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[234] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[233] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[232] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[231] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[230] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[229] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[228] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[227] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[226] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[225] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[224] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[223] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[222] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[221] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[220] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[219] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[218] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[217] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[216] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[215] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[214] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[213] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[212] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[211] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[210] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[209] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[208] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[207] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[206] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[205] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[204] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[203] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[202] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[201] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[200] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[199] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[198] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[197] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[196] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[195] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[194] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[193] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[192] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[191] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[190] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[189] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[188] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[187] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[186] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[185] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[184] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[183] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[182] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[181] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[180] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[179] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[178] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[177] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[176] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[175] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[174] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[173] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[172] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[171] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[170] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[169] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[168] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[167] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[166] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[165] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[164] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[163] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[162] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[161] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[160] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[159] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[158] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[157] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[156] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[155] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[154] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[153] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[152] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[151] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[150] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[149] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[148] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[147] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[146] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[145] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[144] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[143] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[142] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[141] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[140] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[139] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[138] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[137] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[136] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[135] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[134] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[133] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[132] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[131] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[130] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[129] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[128] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[127] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[126] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[125] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[124] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[123] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[122] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[121] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[120] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[119] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[118] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[117] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[116] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[115] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[114] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[113] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[112] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[111] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[110] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[109] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[108] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[107] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[106] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[105] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[104] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[103] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[102] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[101] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[100] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[99] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[98] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[97] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[96] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[95] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[94] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[93] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[92] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[91] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[90] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[89] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[88] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[87] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[86] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[85] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[84] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[83] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[82] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[81] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[80] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[79] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[78] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[77] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[76] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[75] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[74] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[73] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[72] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[71] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[70] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[69] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[68] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[67] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[66] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[65] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[64] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[63] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[62] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[61] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[60] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[59] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[58] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[57] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[56] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[55] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[54] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[53] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[52] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[51] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[50] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[49] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[48] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[47] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[46] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[45] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[44] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[43] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[42] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[41] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[40] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[39] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[38] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[37] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[36] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[35] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[34] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[33] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[32] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[31] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[30] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[29] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[28] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[27] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[26] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[25] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[24] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[23] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[22] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[21] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[20] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[19] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[18] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[17] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[16] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[15] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[14] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[13] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[12] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[11] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[10] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[9] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[8] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[7] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[6] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[5] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[4] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[3] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[2] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[1] ,\mux_top_inst/algorithm_top_inst/buffer_line/din[0] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[6] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[5] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[4] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[3] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[2] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[1] ,\mux_top_inst/algorithm_top_inst/buffer_line/adb[0] ,\mux_top_inst/algorithm_top_inst/syn_off0_vs ,\mux_top_inst/algorithm_top_inst/coms0_wr_area ,\mux_top_inst/algorithm_top_inst/coms1_wr_area ,\mux_top_inst/algorithm_top_inst/coms2_wr_area ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_q.req ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.finish ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.ack ,\mux_top_inst/algorithm_top_inst/usr_ddr3_wr_p.data_req ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_q.req ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.ack ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.dv ,\mux_top_inst/algorithm_top_inst/usr_ddr3_rd_p.finish ,\mux_top_inst/algorithm_top_inst/cs_r1 ,\mux_top_inst/algorithm_top_inst/cs_r2 ,\mux_top_inst/algorithm_top_inst/cs_rise ,\mux_top_inst/algorithm_top_inst/ram_rd_en ,\mux_top_inst/algorithm_top_inst/ram_wr_en ,\mux_top_inst/algorithm_top_inst/buffer_line/clka ,\mux_top_inst/algorithm_top_inst/buffer_line/cea ,\mux_top_inst/algorithm_top_inst/buffer_line/clkb ,\mux_top_inst/algorithm_top_inst/buffer_line/ceb ,\mux_top_inst/algorithm_top_inst/buffer_line/oce ,\mux_top_inst/algorithm_top_inst/buffer_line/reset }),
    .clk_i(\mux_top_inst/hdmi_rd_inst/ddr_clk )
);

endmodule
