--
--Written by GowinSynthesis
--Tool Version "V1.9.12 (64-bit)"
--Sat Nov  1 17:54:22 2025

--Source file index table:
--file0 "\D:/FPGA/03-outsourced proj/05-panoramic_camera/cam2dvi_no_buffer/src/fifo_top/temp/FIFO/fifo_define.v"
--file1 "\D:/FPGA/03-outsourced proj/05-panoramic_camera/cam2dvi_no_buffer/src/fifo_top/temp/FIFO/fifo_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FIFO/data/edc.v"
--file3 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FIFO/data/fifo.v"
--file4 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FIFO/data/fifo_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
rxHwfTvBw63R1D9vcdifhe8htvHmMImvSURzUWZ3+023YnPbcUZaSkQvLy/HS4coVhyHd/mefN25
J1ud7SUWoOeYMaWW4PoNq4GdBNldMufKXEofvOaUpWRRtdcVFxXaieqcuoWbdrtK/+PE5EZwE22f
Re/v/2ZF9Nj3lgcZiLrr2ss1RF0nX69hd07jHb1ObO+660VFrisYwRPvG/CQgAnxg0jEZ8FXiWae
kJFGvIYZy2zjm6gjqKb3TgpN4/WZz/plttCEtxkgj6p74VD7gFUF93h3ZkyzX3275Y+EtukLEIih
wqOxyxC1lToUjmlCV0h/hJSj368TeukKKiHmvg==

`protect encoding=(enctype="base64", line_length=76, bytes=102400)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
ET+2einZgJeeUszL+Z0UulsYcQvlY145EbUwqjYqbEDbqcxIWGwLxDD2IN4S2lNlF5xpQsBT8upg
z6a96OS5JxkEaMCZx1LwMg2sPGCXYQ/hFwP75m8pD9Spw4I5ShpLK+qje8SjoyYGCEA2n55iopz4
pxHyL3kO8gy2nABs8pNlRbEzRHZwz19jpeDjhxpTmTWI6c37KjufFnIvphdQFZtB0KoOuS9Joh1M
xehtKkF90gihI6ud3vazWWqUAuFsNMu7R1AtIVSXdH9nYTYpAqMDiYDIh5D8qwAq4HvEI8a/g113
d9w/LY3AYF7TrO8+8ErqJN753C5IfS5yTm2bhnBrX8Lsg7Hxz7YCMuIApQzyEI8ejDjZHdzQPj1C
xVsD7yd4wNeC+d25i82WCZrrTmdGtMxAftUFJYdGKdiT/UtGs+kG/Kd+xG6dvqJ9oBHHuqNZoiVl
CAHF7d00qgNb0dwoEgif3Xa1NXU7sse/68rwVtV/2BzVafwP9l8TFr/jLYLPPKFVRrPy7bILRguL
c0yT/ziTYzz5Lu3qxHCudJh1gi4jS4LFcCOm9MI0NZ+Zz9mb5FXihmVdXOEC2pPJ7oHx86mnbjqP
lOZifpkRRdeOQ3zQ+SCldiFECPT5d+dLpmI6V1P8XEhRcc+JH7Wn9GSC2gU5TFii/MeQza70fa2r
G7Zd5fe51Nh3VM91/oVfewDWay/NwtOP5jwa3TRuUKy/YbReVAkSiepbdepau3deNT1CWbaRNKam
QHlwZRwIWZ7c921Mz3T/xscFuBe60vGQXN0UVtavs7CVvh+YwVaOzWrGuIa1jiASbdU0/HPkYYds
3tnmpdjcw3h4Tgp/KZBmXJRNOAvyVIh+9WSn/Te7SMOcwOsCcvZxFmArOgyu2yGWIkgqmjkVENUY
X+d8Ze6QxLSOr+XgLE9Xj/kBGq7wTVuuxkq/mynAnfluyL2iPBozDYU4QMR0Wliiy4EvoDyiVN5h
m+W7wFA4+kB3K9AD4mRpaDwNSrmg4fISSsuYBZ0tm5tPkeofjJBzThTbx/tuPBj8ElUjEE4iyPey
4l8hhPRSLQfLu1uIQb8nmkZ3/1f49rpvsFeDBAxhUuo7h+kNpuloK9iO9nJva4bqsqIHEv13PAxs
wP/XFnGOn7KiKCsF8HQQA/orxgnBDutk/M3XfFqqVirJDue6yX2TY4aq4448qoR81HXNKgttQLUB
+mc0kBF/bIsRJYPEMV4sf8y9sCn87j3OL0BCnYeFNdbsDda7eQESaMY/Ixo0O2qD0flhNvta/hlN
lE996sREXdQzzHDZEtRj6B8V8IX3p6U/wx1flT0BpBW9RRzrksTn36qZ+ijJ1mn2DUf9nKN5GKOx
yBjw7l5/X7TD3IaTbjAYdq7NqSAVMKUcCpllpsckYnSOAsg6z8vgKrZuMzBK76CjICRbPbVfhsq0
qNKpCNfZJg/OnTmwK2+faWBRWwo1sif+ln3NV0Ncv840T20f2KSl/8gAg8yy3GqCVpwA4yqVYrvX
ksX7LmJlRWMGrp2z6YzgDSr6pkXMkLcfeGUyg4XtI31J/3X6fuzXZRKdg7uVfXJtT47ORTmwr8d9
E8Av9CNDSG16JDNJ0KjCZU3Q3lzctmqNTFID732+a1YS8T8IZVfRqSP5+IvPgFEJ5g4W/TQQfDLv
0c0Jn8FN9VkKzxT+OBUlGBXtlD9UDobnffGa2udOeEly0aycLcLu7v5GFEotLG1zxQ3q1qyreKjK
947SpJlAXKi236ABKQYzO6OPFPnKjywaB11xscDLhixY8gkuOEHZHoU64Cl4XjGx7jOAcPk5TpTl
UNGJ4CrPl2ucKjBsiur+zOG3yn/GnrhXy9LWRz5GWLJ2KsCoGyETNS2cm8ysbf4NRSu+DHWrWuDZ
10VrdSoKTl+E8NPOEeJ1jYKE3UlR6WdzX9hIckdn8935Vlj7EJK4F3KyEoft8hhTKYYjLtkRLbu0
6zYqomta5+SyjsBhMor3I00sMpoHx3wRKjFXpFt/5f97BqeSl9CXJdMlt2nCobw16X79J3O+Gf31
VtXUAwWXK64ctrtTAMzmWv+0nAD2aRKlxcJkz4B/w8dUng0Us03Om7KUV4awRK0cWZatKVt/J4wZ
FthM1wKBabrAgcHXUbTElF9vUnHWKTT2zWPk10+JArRgboo9/A7ewC1uyPOe40sXLF+bH2KMZ8Lo
Mzv8rI3KnKsveTkEYmXBfo4KReNbjJUmALf2cEG/WO2pO8f6RLpf+7hBQuyBG7VwgGInmvQtR7eO
SC1O0hlH3U8f07t/hzPpx7VPLbDbYNfXE2I51qjPvk3Ic/RExh6tKLy4PL8HQy5nqcAX950rmSds
LqujXh8yvJ4wb2qyzcou9ocB5bnDctM/l6+fkr6YnRDP597J++0IvgYkoHbf76TagH5ckPcIjd36
XcMwT2g7Vko8yQiTRD7ODkJxYsLGnevSgfC8va3odoZTfKyK4cYANc7HDFvmXrrhqy13WLH2ViYj
FqcDWDGLnaOHHfEqJGfuylpjzujnvuCwEQnW2d3RiEtr3W4z/JngGpW7P94eRKHvSiuf9JpfJi54
EI72rTHHGTe6ibUM05aw+iXGNCk3XL8Y5M+YV/M6ZhR28jlSLQo+lXk5905rcQK3ZBD+AhvtljD1
0RTQ5EnvH9wOws5Rh0k2sY2s8ce8qlsE/2Yn9o1Z5xeFBCH6LUwRUsKOl8GKSKOSWQN5Agndghjg
tVIen7/s2VU5Co/cvRJreXOdgg8YEDOI6BZfhi9cxGS8X0BF3kbEPmF13r74KH2v92QUYGiOITzo
iib/T/u+Ehat9gLU0B1O9YCR2oCqdHuweiBJfyVbmSbQ1plekiYmcMxKlx33XRDCq+wJyjkOV8pT
qR+NZGbrz9rc+XUfxhM34PHcN1NO45f9Qzv9NJvRaFAjq/TVwa9Msh/UkLNxxz+bUZBJyj/1HwoO
0HsLRZcttoJOWgceiaJr1Zr1e+4YqO0z6gPYozDnMxiDAA5MmrAOO7cXDhen1DWC8N3DVcCGTXVp
qBA2/40ScJ3myidFi1mE5raJQOylnqzFzEMR7WUoENUV8oGhDaZzEkbRr3OuEIypmCLuDISv9kHm
7kNEtTM1fU0ckzctr076VyZE1s0LW4WNuAkjyUV8HQVNxUgV5dONraWPJqpei3LLmK3OfwHL+pcP
6BDtb+cQ3c55HfxmYpdmN4z3hahKJBxTx3p5bEdPWBDAcehQPr1BPiVqU8ZV4ZQpYw6szVqlPyeE
81GUQeoN7D3tS2MKElcGyGz2sEsaFkrru0laruTi9aK8GtNSTCjR/B96eN8BUvpkGV6GbL4QoER8
ugwAWJ8jdNwF2LafRsWEeEg5es1gWm9hcuGu+P1gEfZwZcg+XYBnr/ah9M0GECxgZ2cdv1uNxITJ
xFzKDNt4wTXvcXTCh6iVgdfuF8dkrG1pM/+sv7uv7Je1ENHmMT4KbgYgaaKI119dPi2y4+rKNbPI
o0xdUycn16AG+23TSRCWNm8D77A3nHuKAO17pWSdp/CfsWDw9Jt1qVyvkpMgxIg6zIYiHv6CbxAb
7SmnoyiqrGIeMuAg/Y4NJGG2kB0eNJDDfBmCIMChqjwZsspiSP8z1a9gGUqlfDCCwcJ57r1EECh2
UVNvwY5w5kWcBOmM/EUb2885lEuofMMniSGsxaVvy67i1KPvfYejmf/qjJ+iKAzPwjPabyqFuFW1
o2MDjctGHWX8iRcVRsN7dW4cuul0QKOY81UQVcVeOU7/bfegabYwTn6Ed6k/ttgCejzQeEV0cSnK
m/tdrGOIUYjGhzpY/X1XKhNR5lo0LbxKhB0ECvR5eMj+MaLV0VgHQ4dK3Ag9t96EWIeAzyRf5H9J
x+Hwomo/ygtlJLEFiZFydOm5U7QCXdtiZkc0IQhXZQRmYTr8arybPkbFw4fQLu2LmQggTv47wq4k
jjDrcWDPbtNK/DMd/D+ErK34tNZibq6kaMLJ7Vk4Vx09QFKmHEHCL7NhBZnRCWTPOUMtuU0PmgBL
CEWWxuRPdZbgcqGSUN2Mz0kFwZVF5KIYL+k9GDBErM/LK8aORacvPNlWEOCOSQ9bUSXhQckdSQDP
jHkjYe2H9e384D0EBR7d0tsICCer+AW+bJZATjYH6CThsgQzn9QQAR8uwZ/eyCQbKfNPJuAwKHCJ
1yDAjq5KQ0ZZGQoi4oqxXtYrI02bpV46xFhT8wet6r+1UfAed50iAsFLgmQZLCJzmaCn5FtTJuGq
a0Ysi1lbj2Kxu2bm3tVPR/YgP2y/+J5quQuvimyp7LielXp3YXDKZ0TucQTWiNGllswOA4v9Gz+H
yyFwQPc29R4qtAsagUWqzMNZFw5yJhRhw6/Pw9MRrNAZzwar6YPPg2sMhuwFBrQNQmFqyMBloFwc
WGvt+D5H0mf7gX9/3M3lQsMg/mutqynbVnxguiiOs75x5j7gR3I1J/f5pzTQlOyM4qyKYW537v82
2PtgVQF4VJlFsemeSr7Xvn0+5xsp4iPpNNEviWqAQYCaAawuSOGqWJ9sRLN4kMCS2p5pHQpdZqD2
T2KJ7N6hMj1RRvib6F3+3hpgBiNgwVn63iC2pbz6PAviaFCBQnbYsAF5QaArJMed9V260mA2o22B
YDmjMl46Y4cIp7BGzFTYPl7d+YpVnRkiwLvMB3LDSLRXmqPNw8IDK7ErDHQcy+i0id2K4rbPLL71
8lbFOKrs0jXNAl9TXXKw6tbQUEJSfGJ0YWIgYcVVnCw4tcn85UduwZnscenYNtksAN9VH2+YJ0/3
fFgnC5uHUjTk75l8Kcne2kDSzPOd57E/7I4U/id1YqhP9VWEO3mcqxg86JX8MD/o4Xj1qCFF42ny
j434vYt75wAe37g6eWfQ5foOqEffEjXkPz1QrUeEDEPAg/AW9MeykSDeGKxzefDVEHf5XvAn6aYr
hzfNH25ORZ4hqa9rAQ8m8Draa208JdhLaiYK3gNQ6ynWcUB+zSYL0nOumg/IjRikdFrrQZNbZI5E
oXhzpdlUXjOsgoDQJo45ujZpJEsflnoDk9fUuZ6uJi5CUYr8jNtOKxxfAd6E8Qw2bY9a51oAbItQ
rk4f59ESDa/xNmrwtF4nmYhNjSPg3I0CWtPnuIZDhOz9CIX+c+vlW3/jFLP92ARz3VnGl0O2YG9B
wqqqq2o6yF6+VfWrUKv9symBTvS7KpazEm96ZrpJ+A+YC6huEz+504YjI0Dtuy344hkUMIMYnocb
03OJSJSFOw0DLbkdWkNeVqXahw6MYwEnJ/CKE5Pes2WDQz3Yjuk9SI/MceVEvAXZRdR03cI8cMRh
L8rQdKzFtd5ZPq34fwDUdk5hq8TrW4iT/mKK3K8yUB9n4XiO25pX+PiCNQRJgbEJPpzVvwBIUk7q
s7+gA3NUpG7RT3qnENKhn1O6rD2A8V7Lad84WLdw9m4d6JD9Xl9WY1B/o/SDM1HmiL2Xg/mxB//T
Q5Y/qNsDH6DSTxIrsXWfVNSUU+hZFyF3wcuLo2CVmhv5TnqdMRGoyG5scZkjtXba4MjGpilb0IQK
HcdedANegmbCTJocj9xIjPvNGbZOVoOHUyUNDjKkGIiyc0pzWkJKRNABewJ7F9NbuVmalDFfRH2B
PlAPiMySr7lwCr0MHBiC3LgItoUsuaeHythjEIBvEWgxRxrFTAsoIq8GeX2vPbTORvux284aGPGn
uTn+OKV9wG4yqWZzH5CEOOIHQqO3wm0wz9KjH68nVsUHw3DQYkfB+ZNEt/itICu5zEfm673IUWDb
XfKY5X4BtXE+/nVIXshuFMCjxZwCI+zkLD3UlkXWh57b6P5sZ9Qu3dRzy6eehu6/J6P1JO2UlAKL
BQUnrledA7UQ8Eyc8oe3XK8ctOURgYSZGiFGnSAw6qxIMAh4dpUT3m0u0bqjFvX+J2AlS48WmMwh
CTjxwF96VC1j5T5Th/ueD0mCDRnnOk/ZlWQ3Fu+W2V+Uefj7Zj8PZqOeTo0nmVmjbuta9finov9J
XH4a7CqUrRgK0mKjQF7CuKW7zKIGMAT+tiA2PEX+b9C/xbWqb2dN4Mqz72FeMBQYsS5D2n+by1QB
IpR4wOVDuOSKkJAfpMFB7YzF7hwSe1mROEQaNi318nGYwRSqe7bvIrt9yJXoYFlAFDqY5/lOHTQY
SIAZoVneNqUmAZpD/EWVMRueJevsNRGm6aLtZn+08OY5TQvGt074ivMy8mcaQHg+s4otYqBMwjdD
BqGcQj3V8YupeN9yJRbNwl8dxAHiNjns9oqmHSIJlD2QTJxYhz1BSSoR4ADHpDpK455GVuySUqg9
3N8lWnrX5QFGQFPBsvFbWfRXtp/9cSVz4uGQ/ydNW5jwWLM2vxBRWi35n+V16V/ozz7/Y1H3Q1N+
IkcW0Y4JcxaJa3L+lpIufQfVm1GsIO1xc6eXeHi30yjRs4ZD4YLQ924FNlmDtayZWWj+PsXgaMI2
mmo5uOh7GNqMYGPmLHZdIW2ivG9dZ0P3YATBZ4smK8vsnmlOwLr8n2C5suj1Fh8iOtbfVtCcVwB+
CuYUx4g9hauyoHc45meD9Tf1YrdafmAD4OiNJwXZgQSBCrFt6VMWyR0WSq3sA79aaOvyWmchQuqo
YlBJZoYRMQNuDHDPu/NOdRTLgPLL5xH3bhf3GGL/za8sdM7N41qkC/oOFdBGWkQMlMAlrvNFai6S
dkIseCj5AVBnvH6lcTJlJGzSZqNzzd5XmKP+iXII72FxGXYbd8g4j9QPzPLNTkVfeIeHOfLw8VS/
SQQ+hgxeUW4zzR0mYkKRh0gng+bq8TK4RhB/AQFcTWim7ZHXdP25nryxZNJGT1zrp+ZOMS7Xd+Kl
Bw8rUFqoOZ1I/EA2Ye89EB3pKJJN1Ebi26liw4tNMOEoPu3eKbLoQ7NYEhT36Iubf+9rCmQlnf+9
w46blEln7Oy0395DCX/UderjbTaNblEeRodf2LY7roLQMyXWjFpg+jk3UbonQ/UX+9GqycZxa94d
wfjzCj3FLs/wHAg6A0nLsl+PxrpnryPVpVOqA1tHej5Mtr5w58iVJnGvIevx/KsTnzU5NRrxzIQR
cMVmS/EiMHaczGgiv3XLB7Pv73ub3v63x2nqaNRXeS/G2Y3UY0AD1580d5f8CeIRk5xfK1u6El8x
vzlqu+vF+YbCD5O/tDfKbmD+3lwpffGhF9QLDm65WEiYHXdzrPhO4AyUXhYhSAWs553fH5fb9aeU
rgmyijZ7+wM4jUVlhUBd8H5wFUCgZEGB9u+5bpRILk6GtBPxa7BpfkPLzhWcYKg2M0p/1L1lJeG3
i527nnzdRRhI3iy51RR3VKyGEPZWcd98WE9fHH6emTOqqrXl0BSicWiTMA5sJlj8VHFCnni6c4F3
K1hG2fVl6J3n9grANr+fEezGJUIF0DZvk+L3QKqQ2Vdu9dzu8YUXEDR468HEqERtYUGNtExVE57x
N1jK7Q3PvIY4f78dzbyuH3Eq4Yf7smiS3RG00Jfsd/PlvYLcZTnXIjx4WtiftgC+aGI8S0wtzzzW
zkZnsXJ2PeCsvfXGYtRbHSricfokvBBM7Pu7sB9fqU7Op9R19KTIU7FycW2up48fRf90cEDrTa5A
qHa/0jVSZ9fe2g5rRz2BNznQ8/JpRkBPfHZxaIktZ0r83LDXqJSfs/X1/U1RMzhfEnsxKD72NZHY
4RhBKZ60iFCra2UjEyA7CfTSjfms0h0pM4NMs44kiJ0E+8ZYZFOCu3BN3rX9jyaODryUb4Jao2kX
uFxhp4VxAH2rLCvT7dFv8p5KvzfCJf1/UEgYlcWXlJ0/PowhvR+OaDQt3VvPQyk2xvG4bL3RmnX7
gvDH37+kc/1sLSm88GarSgGUYTK/Z97lJp3V14erPeNnMRPoVjXHZ4HkBesuG+2ri/9BO3uurbmw
VnLE7VskwRu6yZ98+Q2PFVJkiirqXaOhJCzhEMMe0BYvHyJkzdIskJelDCkPCrFPoCAYw07Jhhxd
EdpyG9K5DGQrhHtlAK9W+iCuwk1hz2WQ+JpQrVfLhdIpqHhrN1ChUCeBgB+hVav5WqU63j0YPRrN
UdjKfjGrwDd7ZTRNTV/3RKuZR7kQ3bJyQow5jyHI4m6bLVJZmjjG3NYpl/vmclS3vj/LX2NnEMzK
8O9CaPibWywhhz4GobOZ8rjnVwE4dO0hlaJ8Uer9/Gy4gIod0mWpfVHKJUVDpQxV5SJuBNCb2oag
NnYuirL5rAK7uRfZKdNAZGvxrFZfnx37Lobb1ZwCopAEJ1VD7sa3y7JaNzzj1F4/km/6HwvFQ0Dj
Acs7vFRmOjWCLYnNWHyxXNyy4w+EbSbfcKdPAJ0VTy9u2r3E0JtfOPk8wePlOOL7UE9LsTE1LZMr
VRng1OAn75VNo/7B1iFFf1oOk2JrKreaL/Cp9g3z7Olir+q9F1isFZxcqQKx98sJlODQtGm8K14N
lEhpdabhwveJwuunyIWmRPh2gi0u7Ngutz2lq4kCJFaQMyploZ/zZD054iNoquymLdwjugJfwc0B
a/K/wLQXYQNpaQisSewC32kqERy1kKWNqVwaFEfkyVRpqTjWWF8z3S4u3xkEjIa1GfccuhOvNqeD
d6/Ag8021P6Mt9NawLbFqGKdW3KyFvNwWQ+1+F/icJMtkGdx1V4+lCi2vJiUzJTYiPFKLW5UgoM/
mtigerZb/g3iLpDf+WHIym0PB1qYVdBG9O5cNniIVWhkCL9tFNNSIwqvstH4qwrc938OXqyw0SFh
ywfuadOhEsqIQMCiEeiRITdaxXQq9cJPba8ceCQcGYEVlNSgFsaPkQVYT4WhWeWwG16mQhSdFZTD
O/9m5ceepKw537sU8MQC71EUofHk7xYC0x/0CbCD7/N4s5lsup7GRfF3zLyRYvoThVmDs/6lKEUw
eKANVvVcP8AApmhNty09CRYTsdqXAmJx4SeIOmxqRGg3m7xYWUKAoYq6MLrNnq7VhqovYxrHaKln
wLI6VX/k9cQhGHBBFmLA+KqyXkiHPl/4+KZ457Th8PehOndkC739KGWSunBoyidKLvjfLBUHnK1V
b07FTRbJrbCoiHppRLaxXGT0zDrvE3YLPslrZIq8L4Fb2NnEcEfVq0DGv/aUv3yDhhLj0Qykik9b
mWF1JpoO9r8HKiOsPB5Kpers4z/oZTPyUh3f+5DuGKkX/1WwJYiDzJf/C9b0U92CoVRP8qn8Ztag
/Ot69YaQpJ4jtBslFL9pwM0VAahYjXGgyCQKaUWnzrdsq6a+XBNxuG8qtjMFwlUHIq4Drjp2sQ17
0Goexwr0o7Ef4Tt7HlpEjccgymvIzq4M+9pM+h6h1mnImZTRqtc5PupFCVY/05MWQT187nBuFKIm
/jZHFN7nuO8xHeWuUh5UNFAaNnrrOE7bECLKTBzJWQIMfVvE7AVfyVLgb6AxItIxULja8/VmV0MJ
DhgJ7rhxxOzaBaGuCnPlh7oi2bFg9IBMylWPCmZnm74Mdoo4qWM1OBtp86iQTwf50W11knnBILDO
i/zI7RMnEI9/htu4E4hGDe+Yofife+r6toVgFATwgR7HuPgFMnN/8C0Mk/qLJLbbsSw4gzFjhEr+
aamFo9ZEcUljrxEW9CyyX0xShT6CuYvx4opelCHirXlFnc64+VH2uiDwvpiFevfqRuyHwvcl7Koa
PHnFYrT4EpZjj4HSRe/TWsgP12TkitYEkLkuP7FDZPgGyyPpDN8Z+Vx1fkkPmBW+RPaDsUadAl64
/b2UV80pzIE1QoPyPe2fqSVppd8km3DN613y04agO0lXxsfhE63fF9Pf+Y7ury61mJMgY1qXzXvG
wrcJGrMAUNz2TEcGXbcqow8R45VP2MztG0oR+FqeMpB6HdetKTTqvY0S/mskoYcCuU4oANLvf8Pm
Ijb79UddDVWSCK5x7nOOjggUN0e4cQRsJbByMUvqmYqcJdIzf7wB/n/hSmy4tpBy1FCctNO66X7k
zYB5BT3L/uV4hNnMjGdNS3zNVpaK0p9oS4XIcZF3nuyfhmmNVtYhOAnSk5LNAt4jHM4TSSfxXUmZ
3JsbMSOFnmKKaSyu1UZcfhp/VhRcyLCCaQVfhdKqJwQdpmyfF9GOheDRiUfg7kPgve86dMHZW1DW
etskNy/kCbqky4ybPfAw6+n7e7QZCzmZ5zAL3oAzj9eoNT+bfLPeBvRiqCBO0d3C9KSdwF3D2sTY
q3bqyzCSV3HLZmRbZbB8PjL5Oh+sltI2D8qnGW5qkUTvRswoGThdPkogVN9TejfTFVrAwAqIp+sZ
nvXE8+kegV6jwezKGHyq15Coz+rEo6bQS1xOaFf8vJjYkz1+mj+KC6X1egk71WsuYBl1w0JgRhXN
Z1fxLBkrjSp0KNYrpGB1nLhQMQuSa6VaQX+kRCkxuFMJGrkMv4fs4EYuTHheRkLFji2mBETflKcE
ncFPWOkTGLogFPMEubq5Tr5k0Rm1a/4xaYz2ALeorsyeTO5AE331mWy2EmH57siI+wpEC8ixoV/W
+hZtjimc9ogYGMiWw9z1L1f6OXJ0MrC6TrU2fS1ka1xkgcvyq0r6wYByBrkAmeI7r+T5M2zj5QfC
cBJdzPG1rQlLx/I/C8Yg+yHn4ObCIEefQqorZWM/tKRnyf/xbfM/rWVJ9SiGIhY3U2RN9CUeOVGT
qRl9bfYAjfKbFv+5uR47Iuvvj8AMkoWv/3ADlEsCLt/0MjblohN75Kb517AhXgvmKRHocHmP/k4n
ynHDSGUgqM2NdaOfcI10oBwzXYYM3/6RsvKKFuZk2ILVZFfsEuMibVCZMmytbGTOuHb9IKrj6nrc
a8BCwt//B5zNZz9tSIHAKfzXapGXYEwxRZi22tjPI+saQKQxrPmM3a1k1Q6g1cSolXWxfJir6oRO
UKQDVNsU48m1QuQ0T98Hpwk2Xzmwip4pFIrEL4+Fz4pfA3IszXV6saGBYsXIZaZnjMvBSAzWh5Dv
b+q9CyqfRHEIPgD/JR++NiPbiRa6QO+ZHdt912kQKNMq+xqLol5DlUse7qC6vnwU9H+J6I8+DWQV
yOoHaVaDH1fYLMeXDbeeCt4UKzOuxk+F//g2qOBH4QUfkaPN0UdXnQUQEXW0k0H+aTOtYUvAVCrR
OgizzVx66CDGVU+WeoPuILDKdA+Zfk7tPY6PUgDpSDMhCUBZvEnZMouWjOr/Uq6s8ii/TEXNK3cy
szDCGJritM8xZDXyFpv0/gZRBaTEKQLaIiHRtFmPkdzJgglfjPoCN0yknNFNwzOx5S9mnNatG8g3
+yvSZsqyvxxVcMNF6CuPZnr5q1ErMxo2KYUTEkx2VnIf7JP5dwNVshM6luzCEHKfpPI/NyIaREmR
Vq6zzxfkNizz7fgqW4/oUzt4eT2Qgh8PNtD9WsLNYTR0W97EdogaIFzT1mcdCX66/S9s3nezbMcq
sibF2Nr+8+3U/HS4nzkqADGbfbzVTl9QX+fL7jPmRbP5bAtYsXV1rg1g9O1ONOEMrGN0ruUUYE1D
iXIkudrpeEzjqEIvkozhp3u4zDWBvhayE9vBpo11fxnvWGENl/VM26d+W6eXopP4mCm5sYwavd8e
w2QMkbRYQ0SovYFr6Entwh/joNmxRvjMUYL47/L7mD7t71A6bZF6csKwmivpSNC7KfatfmWloWKv
bKjeTWfdJSvjNLGhpT9fsLaUWCAypsfrSm2qj7gvLX2k2HIg9hLzzY26JObwqjxIX23k7z+/gg8t
740YSt0tyqa/2cfcTUdOtS05PrVQwspS/tu51v+ZnnGGgQMIC6HdSVEjZeg5zy1ruJgLVvJQHUW1
GsXXu9+hxT5oaIjOZ4o66Lx3XYLD6bAhnwPdQtUYqIFw3C5LlPKfdKhcScdqLgIMuHmv/BlYyZZj
t3duwuaahcDcxwJZ96qUKgPX+eQi3npNH6UDbWu7JmMb4jxfGfcIQczGq1/8zEWbzvibe9C4brcO
JaIyvTZKwZPrlpsf3pPDm/ZoW1iHcaFO/FWnXFk7324Kuz2FTa1ZAGe3Cgn1h7ADYiiZyoR4sTNB
TwszmKasRD4GQg1dvSBvCs9AoZdbYgyh6ZRf+hXYKlcmvK+nzQMO46gm/abQPLhhy26jeACt9J/Y
ld5+GJCxxchf9Bhivm7P1D6NfAAMxC0dlYkxfbeYin/HSVqcHS/kHZEPAKgE6YIkN60t0rTyshPU
po17PD8Nk27O8i/+ai36vEHnyxzgGZJJDj1+ZfWsL1oGJn24paB/yXvPdrs0FbhjhLBhBXEkHHaG
7GD58d8sc9CWW1yUiRPaZVsD+EJ9HhA8uD9Ba4v2LzYHi5BPLFvbyAUBaeSp3J6wqfCl9Ddq0KV3
senKkEXKtOAEupFK64MauWU0ak4/Xxj4s8D0jYaBdA0TMItwHpcj2VxGZTmlu01P938Gwpu92Gi0
sXe1zft0x5Tunjb3R85v/CBxZRwvEShGk2bQJzNgF6ymaoxVrUp5bdaUb26xUw7VnXldj2gT0chu
x0IDGIsxMnV1WdqZCDoWXl3+F+4zUWiRh0lBMSncBWTnbLrECq67Htvm6kG8MX9+KccYjQMVNnv7
qlo+E+WdOk2LE7nl1V3jyd9QzTKSUr3Y9rrzVdGwYMBZSgv78HbYOLNPTER94FtdRfncVy04+UbB
cZcXb7Wf5Kr20KYswX0C5GWuyT8nt7KjyIDXVa/WpERpJJEc9YOUILMbuW+jDtnxDR4f17tsODuN
EnJaX6ZK99aHUR96/d9mRW1NJHr/vTPrQowUqXM98mLr1tCituIFuPAlJTyDKUT4k1OeGTQRTvXF
79McEuEPJ9TBjr9DnZAes2l2kiLeUtHsoWAIBhLZY6AL63mr5A+1fq++C2bt15p9cSPlv52B/cWx
cwhtMYZ0A3yoKLPw9OSI1KuKgSfR15ojvr0NVGhXT4sAuHtgOkBM21l6NN5G1KdAAMF8PXVSxgSi
MpsdV6Lt6vQX9gZzLbOhV4glHy3A7t5DwRPS81R/Vd7R06YFg935RVdh3vVcceAT7g1IFrRUqQse
J7lmiq0RYYibZvSVNVBWIjcmpj9NRHmDZCxS9ST0CqPxZu5VWBwrXzec5Y3aDmLAeCiIjMtdZ5TA
/MTOo10rVY3npUOSwtCaCDXCAJ3QvOyjjqVO9C31SokXqdSyAYoewLrqxWqUXXzqJyec52p9tm0G
sCcWjFF9n7pTKkru1UJccTgYpw93UyyoUIf7lrFdivKvXcrJUW+RmamqQCxMMDw4flk3BVFfelHh
XpgDbCsnMjU19VugqrilbflP+H6NUVG6mY3i5QuxW7COv5hpz6ooU13mM9TVPe4sVfZINIdNdaO1
3iIU1o5IcFl9bk8UX7XJEwJ7zRhCr8VdK060fUXC/YUfNgxX5/hRsjQx8HB1zq0ph39Ku8SfkFjC
cUnlvpVZX2quLStj5SHypnlbESNrrOH0txWLeSHhClCrlVi73khqUygvJeOVTr+FnJ27GldKm+V7
NcmOLXNwGFjYbD0cZHY3qJNxy1K/vnc2Caq1vJZIDQXQI8aFWaCF2vRm8DPfjnXmCAp+62yGi9md
qgpOIe3ghJnsjUMe33lYbErM7I0t+5xQPKvOTXykCR/IIYvYS++j/4Oqh3KXNo4h6BZTLogg7ln4
nGSJVi0OPt8q+OOPrPrpZGa6v33zEG3jiaTALGEUJhiOpxY1JGnFUSrE4MqUcuZ64dxDp7BNW3Ci
VWcqdni1PReETgormCWG6hX0SVOywPqpu2qj/uxpBgqR6Ma1u12q3D2FyhNj6d+CL7Hw/Eai/qsB
1vu3qyksCUZXFeKip5BU2O3h3N5xtItVl1nO7YM4ri2eA4ayFExDklRVchBqRp5XCxmmCeJ9sytR
60/F1bvxhWP4kMZdgEZPTLRdMO4adFL913Di5rdD4OjE8cRRBHv9j8IcuFT/HzIbfB1iHJgEjvap
uTYTuFhedw7aDAiHqNaO1zy6vPd9gcmVTCcIFfwWlWJ5ukK/MRKIZOZY9AfQ4Cz3FsLXIFgNNnNS
AgpgyNLdSU41/Dg8RH4jRYzOol3L5vFexiqASYxJ7w2PPUNtLew1GkVD/6VQW6BShMBLzkeZEbiF
LbtQKQI7EnBZGRLIfNgM70QO6Et8uO4feLPY+SHSn/kjxWM3rUHH/kba7kIDZ8AlomKtBEOI72EK
bTJypasXLC2jTkqIYZ1GhUciioC1XJEIYVIpWIZLLwg/4WPYxxmERHJKjiMlCLjdC3cCEoPEzEZd
cRFrdu4jJdgaqMUfMcma/Obkn6QiI8hs4hWvXa36tkQgbblCzxoiJEL8R09Ok9/MD1FhI1fAbKo2
dfyrVzMl6uydBszoJqpXeDnrvKFIiOkW59o1ZCeg+Slbr7XjtYhXYDsnxBvJlRpNQWHzOQdH5DJm
oteffFG4DlqoKQPidt4idV5RiXpiZ6Ox/Rbesj6lSC2iT2YW0ztA0kpXVerTQU4TfBf5Ko2Ksm+T
Nd5O3Lr4wvPXvIUO8onzpU1Wd7GDH13MzcN8jLhJLqLDJ1kHKiHKr1xKk/wfyE5RjrtEoj58uzTq
AmgpccDzzpaL2ww2vLsviIOxZiDx653zuBT+ma58QkUfpcSwbZuPH1ARLQgX0Sr6dgOlyoEFCuLZ
L8G1MRZlLGjB7Gh+y42o6KUPh5PuJzcMVAZMPzmjC32vkpLxHeQ9eeHiWskok5QrHMlgGDpQeopi
xRyHMlxaxxzGs9wotZAuVuXTKhcHFlcPNDdJagTxb2v4Qrf1K7/WIANJ3hDyzY6fJe9d7rxgvcWX
8wz5ELUydRMkIBRCcKIrjIlPFE9kEE5uvvEBGEA79AKi+5VL2I5xTXMuL8DrbMRnce7bUGw96Po5
UDjZGBoht09d/odDd48eeJlKHmiOX85CRE4ir44Tug6z5KnVgXIqZr+eTPbjsSx4vOIftDSUVchK
9KQ0pEdxPTtAEtzQ8CjJLHkXXKORkoBvRywV664EAWdvg2FhmMFQ0XDWCqmVMLQfdyFLzg5sYnZH
TTYpDN0pfJ8VBFjZlCN/E/GIYC40VC7uzECjdBeZXa5DeMF0Xxzi7GsLFJ6M/1xb9sWBjhHAFhh/
Vmia8mbJtHWbWM+WfoNMusF+O4rJGw/KnPYXKnVO1E+cE6Y+DQrqJy9cU3alkG2APqc5Mll9KMwN
ymT/u6EpiE2CWMRmzRc9wtGyF3aqudEqq2B+P1NEmZ+DPmDqrIX7GDad+3KNtL9ciISjFBYV037s
TncLX4HjIPWsm41Kr1d7sjLJFn/wCtzAJyDj/p8BQLHl4gcgXzIj/FdwuiDXZ/GOlwGLauMjHCF5
o9x2yKnn+KmUHtAC+OY6+yqJf0OAGTCRyuCVxgrSzPOGipcsCcKirrZ8h9+z/wt/YqOFxw7sCnIC
qWpE+oHa2XJdafetEA48GhVO3rbTC60qdUVD6301+ls83vpOcch9/0uxRQniSnWE381dn56y1+tK
dcj4LGx42u8IG0mSQGflblmBXV6OaPWO1+KIwJyg9Co3b05tYtAplYbdo3ghEyrErsbZTbl9Zj85
uOhz4RdE876BNRrrRIsQyxbQ/HuJ0J0rOhTggbdV1wg6lB9fbQlr449MdPhka7ZxbecLF/zqCa2B
ndi7mzZgOA+5x0qRbpEFvb5ZIaxdSs5ooLYLCWeGJZjquaUBdcBubomntH7dp4sQ5MRXhv3D7+OZ
YHXYwWW2Ak26pE5kvNzA5A1CK6c7OIgipRLaIa190TH4KhwZoJI2HtDv7Jfq+gOB0Dd45hMSyr/7
avUvZRcKH8DV5m31kuwZIkaiTc4u++yezrJEzPq9T/4nvkeS7mLyFLInTo2dweGIOvxfc9aZK64G
sntRbMXnan9wuJeOk4FPMzefkOc+7n6GZx1PX4ufE9ZYrUJNeS3N3JNU15LOu1OQrT/IhLRLXA2t
qm1Ue66G0CwxeKNZMk3Src1ob3CsQHer2oOp8mZgbGAEOITeWUKupP0WNPptVlI64hkhnFd7A9v/
CP84aG6LbEfolQFtmN+zV1zdwDkSU6z2xWH4uA0DCERzUX2XebWNP/VZS6qmttNxBsDg5a7KnqcI
vak0KmkCEv7m8vXC25zyy7cAn++1CW5rZAtAtPYGouMVNphV3vHQ2BIgF9YcMUsw+kZIAR+liCNC
PTkB1SsI6a5/k30TAqBBl8qk7RkSAsWOxYrzgrQ6uOXPrhb8957ZMf6QkG37BxKwgMxd2NquRVnm
hk8qsSPia2i9P8C6krs17Md4ZRTOsls1ADj6rTG+hzndaBw9+MlXUqmrdyu8ip2iR2s/wpk3kG0K
i5PXldxnd5HSvG6orTa2hTAHozcOTa8Iam0rCB4oggpiurbY3V5d09NWag2ruVWotR1HkPVXk5Jm
d+gSYnmxRtU4/C55MajXo72r4PI56tyQG67o+a2Epix2LNCEHBRgaNjWM8a0uLSN2NxMbpNs+iAN
/bV9bAxXaflq0DdiCLGZo6aVu2TUjzddF3tzPb2Gr0wFWVxwyC1wDxsou43GM1Q6gmRacr+Obkuk
+SWkQuEz/MQzdsqsgUYlQ98SYojRGB1Ar2/wncL4aZCD5y+ZUyMb/BWja24J3g7HLUv4DuWRJimg
dHvAR2+ja7l3NBhDOo/WaFm5s8uz2UNXM1qwUtYNw+xb67sadfIbmr0HnyH64En4gjrJR14Zyb4X
Bt+qFMNk6IqfTXmJQ6hpRB4c7GjO7ndjh86MJTLX5G4xoDSErtXFsiYQvnpbqVAI1r9BTIvhpHov
cW8MRF41WVwh9KFPMwsKNbXBIQVeYhdWczhOxoMb4vFFm/MYs+UxTz1g2qxOyWf86iK0Up7J1eVo
GCQuTyB+jStVFi5I3yRrABTQ6uQbk6+f9MZvfDlI+SbXydo313vNOE0Md1SDwhvW0ugpsBDy4IvM
5JBfPcZzaVGKl5XS4WyufCR6mEEWAJao9RwqxHNuqaXmMqnjryY9FObrXb7+/MuZV9J2euNrjC39
Zn2KHZza+uhaESPamoW9gUbvhTfF9Hm9SX9/qdqwDOlovqeH2KIIIIGejcKfjbkMzaOwDF0ff+eM
ep5To+PjR1N06PeGY4eImoIX4Af6o2IpCEWyaZLmtJ9JkFbfnl5xGj3ZrxE4y+WsKkA3239ByF4c
Ooo0ZkyVetdmnTiHVdHR5UltlU63D27IAPU8eV9UQxqV4gmMEVD6cN6Fhx+UH/OBUk/RAqzidPGA
m30PNU31vkrZ3oA1I4YoFCkJVi6EObE0YSUyA3PBjMvSIeNSrA0F25v2h9Vbvi9tYLuI5bW8sSCB
NR5oTA2iXHcWenDufER/bJy3b01LnF6PI+XF0mgDD7YTXZsZlG29C6fuB9dJpNPYiQVnhYNET5Ok
iKGrbguyNfjoptb+Jh8PcDp17NzzXF1qJyjW57F0Q5CWJVfTD8uQ+YZsWQam6zn07iXfR87nptLP
YuQRaHf5tK00NvVZ8H+3VArG66JV6ieZI9QmtUs8k7GUB3kqZ1qsDkxxLkmqjGQtk2N3Tkjr+hf8
6vId+nlh8TUq8U0ye//30ocVfuqzrxOhTkI3O/+wSTO2d5sZ6+5r6U1g4LgblW/KimmN3hwg/e5x
H8P+exBZY+2MFnjrtFn3WAfHDIMhezCyqszW/avRHcv+CQSSw75yhGrUFcBGBdBG0NbxAJFy0Tu7
MoIQ6Bx/d1KEUldgq27quv/UHvaiVMvVKR2DqhRn26EBE/1xSa+pJzggZbeIGQAF60SOyo+DKw1t
7AsSQjHPPjB5Sdo77zqfq+7M0FVDI3XjJKOBa61iNcBdqR4u98CVdL9FCrtXN15W3niIEMMbVBS5
RpEG/6hS3hdgDtCJflp9ZD7xDbIKBGJ5aVmrVCPRzcSNK2hNkPrtDFe8RF4uYRMpPDOmZu9iP8uJ
/lglLbi4vT0DuScPLZjNrf00tp/Li8Q6hSCtEtZVZ+9cXPr8JSP4dNE4vwwwLIwRlUcWfsc2aurl
hIRF/+SYHGAG1vV2TN4Eg7uo8IcDP7+0dAxnvM/t2vLbZopDTsLgu2tNDxdqdqvBztyzlly7k5bT
Nu3h9qtdp7p9KsrKC3bz8y9RW/QYqz0B8tLQ2ROZCdpi2SQgrJ4nZ/JYV56vEmi5HunTzEzXw1QE
hEqPEDxtlJmDrsP6JB8UI/ykkLXMrR0KMHbcv5TEkZY13WzIlc7srgjhbzuaiYAeB/kXMgA5fnb8
PztbplGPnBGP7D4Lb09TFANt+TZkSOytHXJDOT+KJFYkcEoZ/eS035sa3COF998hVrCoiSGjeKZc
YoIU4V0pkCSqv/1Qp19XEvwxWylcF/ray8Eu8HbERxUbPzEyjF0I2M0fT+0IB+AxekQVR3FeFgsB
ABm1iHVwCqBmYlKztnKhO7xDgstd6XdRw2qn7gnt9iOzjBboI/3lCaRqWvMeh/SW4yX8FkdVaNiy
zdUqah1sK1xXTzo87nCONX1ngjXndjEEhKUz4wa/v4IyyLIyqYifbDj60hAel7lDSId4gCShMh9g
PJwb7BD3xmcMr4Dzrd0W6LsTeG5RZwWMDc6R0oRjH6NT6/d93rha574VdRsHLInTT95Z/IUoN3Lp
zWwxRq6TjAwqQOhfTo25QChcls7N8mS9NCixZSiUlvSKfba6ouWB28USPusyL7qAj+Pi+SuBL0+Y
+mbM3VWeJsgQmMwDw+iXVq9A6wUTtiOxlWh9pIQX9rQ4dlgfWloaAWy2H6ks+5zoz36KyOzFqZae
AZsaw3aiKCSb2oSj/VI0ZUsd0z/blwvMdW1NpEx4nstaXte7WC4K0z1Vqb1itW9i+j6uZHjLveha
2+rSq7nxiZrgpvZnqDteAJfTrhxyu2E/Jvsm4PIcQPYLosyztwbuuodtVk+3FU4kpilioQnagVx7
P2gUi8ngCi5Oj6voJKazXW0p2SIXz0SJSxq6wl/X8VnhT1g04aog2J3X8+uXApCpHQ5/N54kSz0S
O5EJDlRzgsunOHtXFaNzbYDwXjcePli/0lcBL8qICxsbntgcswZIvMaKnhjO/b5v7b7BToJ1vsfR
cyJV/6NQzXRv41a96y3p/xuAZsPDVg8IwcZWhHO5p8jmVfNuEZbVlaf4ZcKUcuP2trFIt+lh4oOw
bLx9jbVY+1K7MbFa2UbSrrl9mardTs8prDR1NEjWnCZTFC1jYJrmbMx0QrFSEHIZov5G907nnqKj
cOmnQEPqoKrsyUpvvi8zcTjq14znukMiHqy85CAQY7P0w8esSKtzzUkR3IfZKa74gLw+hLE+PBrb
wOYFOGSkZdyBsarUiidCyFN95qam/HoMoC/JR356VA9i8RkC3Af5RrU/UUq4HCg1hiz6USG8viXW
xBY+xSlZtKEb9ntJ0C7mdk4V41Udm6MH2vdEWXPzqg2FKNsPklrPeh5F7pBH3oJHAoy2VnqxOFss
iKLU2zY2VNI2N78wzOXhKPL8fpCb4myp6TCE28EFEUz9VK20xTeqaJMwXIoSFy318/L8ipJwRFNJ
DjvSyowlork1vbdPCbX3hXmh5EhwihnY2NJNpQXPVyi9bhnqOaFygc3a77FVusg7EeeKItmUW34u
h+KaINqFEFwYu2LNJDbBiCadVfYChcFFVXWKtZLBNyT/ZyBnhg1ci1TYEETh0BLe72rElts/Pfdr
u2ggdd49Gi2rhZGaRBr5LEtgIx9vYNsUHy9iYUu27WmMpO4s6fP0DHs3XvaX4r/pQENPD70aunJM
ZFTeJcX5+Rlfafk90IoH6mwR8HY6aJg4FylKpb0Hms3Ubi3j4bQE4ERjezGxs4HbRCfQYHz4881o
sxXaBMWB56aYYnAmNzFyvdqzM1/trGjb/hkg/bVN0bYm1/BPRSGM1XqKuaQJa/VOpc0Yc3T9Jnmd
n2HZxYTQ71d0BEpF+p04NcwdLj0xC+PoXphqfXRV+1QtDPZW7hVM0+tyJS7XG9sJkiKvTJZ8mQT7
1aYOaiqsnxP5Vc9wXcv6LYaZpHE+96eCIfG/ZXArgYrvtH4Ramec1Ep4vgfHEXMgDIivcCeaHP0G
iTvFTvOvUjQ/BO5mpoB1Qr/iGeZWzOdZeL1iiIvI7iFaVVCkij+TFF23xS2zgIGUt/KfBpfnbOFK
GVB3YRQOU5E9Cs4iX/LhpToct9bW10xlIpn4SMCoA8frJXxhZVbHcqMrzfcOpH7WZVFbjN6j4YNv
c4EjK0GPAlGacGli6zl4S4r34qMbBpkCqSmKHsyupMmt2mPFImDdrwoDXfT8se6tLH4d8IBX0Fks
sA7g+x59AAfw91scP5mXoj87eKQYPKGim6+Nk17yr8eTAF327z8YwDolzjbdrz+Hmf9D8iumbKOL
v5KGpfzWe9prWmsWXIRaad8krY1XJQy4OHs6Tudvd1YZMPrOkGlt9sotIdGFH3EkdH9RzMoxfmQd
ggGGfltwamlV4I54u8PsXivh4PWsmZ2EGgg/v5s+mZFIjttS5ZVIkYMYzZe53rwkglwM7/eEeSXF
Lp9hqyh4U3yKXj5FyC4+w1Zo4lYiN5HATBX1c2nXrXYmMs/KwAYWjKqgZEqD545xIs4kMnyMgL24
bxSVFqC+joiKmjAEwSbDgkubWwWLQr6wbgSsZ56c2f30eJZnkJGxiQKwa97gn/tiQiOcZXWyo8cl
CEpCeDpLr0J0Ov9WoTRUHiAKK1i/xMg3A3JM+gEipOPp7J7I/Skeh9ImhCV5NzKVvM3RzKocWuoQ
Y8TsvYZQAyH+sd8t0t983qIAXu3PNUl9ip0261E6XyjIxVP0vk3+Vm7yb5GRe7eKtT2eD5tuLFYd
k4B0iMIzRQ1YhmKPMoXYtskBzK6KeaBAXP6Y8gDoXgponi2e5AwWt3ujj3FrNsgW1K35HWEVF41W
tsR4yqddq+hjMTFPnbM0UlG1jMqqGu6zJn0KQfQVfIhAlWLEuMcGyjhyE0nbRx5jNai0J4G9tlmq
EH88vtwcKV7d1+9y2fLgXk2bY2CCxITwUjH4q1KF7Li7xQ/hZcK1eGSb4uhzHMSNntjxWu3ZE30K
YSIBUVhhvvHIPAOp1Fu7U2wgFm4KldMZsRoruXcYn2ygzHfHNY1dMwnM0wzR+QNTcAIfXyl8Gbnv
ODkFhjQjXmYO0TB8BXL1P303xGgxmrprzHvG1E12fjDWDkqAy2BOJiPo/+gGWzPcehN4A2jclD0v
DurCXfhgld2LjfMmS2UNnITt1LRkNpTuISaM45zVJXMu2PLxw/dR2/g+F1/nNv46VLhtcftd7k7f
1RRfHzwufG7m7d+Mp2WzYCn9FSd+D7tihlDDxnIjec5z2RIjmrIC8qNG5xhX33ZGBpZAc5MKV7gP
MWNZ+yTe8X6Cc1Vq8XSELZI/Grrm/wT7TS94RvxJKmwGiI63JT2qLfCwBU6vzp7Dg+so90/f3uK0
/rU0y7YsKkkkwhE6wFqPwMFiR8zyItor6yJBxrqhRFni2W/FBWrQP+CZENZyydc57SHGxrIhgagV
5ECRp/KhginFkvPdOZkVxxjiAfk7K3ola2NJdtikwuTsvi/rFAY6A7hEHFAgibCmx0T7YZ+Ndhhe
VoqqSTxOvVVpa7szCf7Du4nNp2r+Zx7S+Iwjej4TlyghaUXWpU3FQlrnIoyW85kMEDAlRHqgG6l0
visr0sXkjmBhQ5Rx85UBbrIOn2paM7JBvoGujpS8nLh0hvLEyi+/VpeFZjKnuf2kEZimJHn433+e
spuTnURVb5ZQq0d7W4XR5y/sTozf1mNDymakaj0ZENdoNYU78IQKeL8cn0W6HNPtxW9bSsEqNOan
pfBH2Vwjey1ve6AH2Uj8NSr33hDUpF+3U8pKw4e0Isrq1haYYol18YME+FdO41hwgEbBMPVL7QK1
ncnld9BB9vs4c9031ue2vrZeaouSRCTar8a5GxLJXc4x2+BASFLhTSpUsntb47cjJu/JlS+NYHPb
0LmrfFLk6V2TtHQIC1zTZPcClk4dkBc1OoMqNCM1pISU2Hiu/PdG2oXcqvzp+eWrHrgsTmjv1Uni
AYBVuBjxSvQVn+5IYA7DrQN545XM+gTpwBnRxMIJqLbHdjhNKsCFpmPA5WN10LZCYAIjYtj72XXp
itosClP1DxLd8bZAooH3g0CpQOvLrDiCoYwgXFunf7OL0a7+UHkx8qtpHmr8hEhwhBpYn1pD16v9
x3p7O9t8Hpdw1tzk7e4WK2ye4sTIZKVdPDankDYRlIM/aLjyIk26206da6AHHyED+5x0YJIwml43
v7O8TODiH2sFGrtKYFYDH9tFVTxR0Fwjs2qkD4Hunjm1P4W8bv2Gj2JpGELdYRHx0XM4uwX2cru5
TK5Ygtqc30+NT3V3PssiVPIDzaUD4xise/kbGYaQ9N5NDFUmBK+FTL3hoND2R9/gYKFdEQCBOKjm
G8S7q4HolyrJ9Ev4nA8ojMG5bwFqHkBoWh1ocrT4Z8vq9xFnSKz38dTNFXhm8RP790fz47FYFDZ+
BG171yeXK6xty4DJyxDBD4z5rHa4pk5pjSiX/zTfkAP7SZQK3Lyjqk/DfIvdm1loU9PgEo01aLAf
DZLrbUUtTFB3GqAzgTUi3ceaXvwgHMmtjHwDUedStLaoG5ZPI8mvtJdlxJZ89tOW+cvjRGvnbMRI
DWXEQ8aFG/YX70u+g+b02ZzqSHm+xaZOBGApf8asxQHdrzP4lcIPLUBbxXe+buf5gboTg5PbaAEK
WXn8DBLL/OIaGeBPfftJzgbBP040UerPGmqrxHK2Cx0fafTTu73HIddb3ZTll0GJwcercalUXSF7
+KgJTtVrxaKvZ52fC7tq4kt3+dTUsbUvR20Kn9BYZHCxGkQz1/7LYrxWB0XPrIrs+LamI/LvtGNW
JLRjPdOG4pIf1yDG1l6kZjc12wQuGIj5zVbAJy0hMPBMka/pK4vqGdkMDUqcIn9aNBFi5AdyTtez
8HNovk0Q5bQWXrLlTl5IJsuR+5S2yYdKNctN3xF0LyGWY8WbNpY+jQuQQNlOtHYh7i5kr47c33oj
lyo33vNx9BVxROPIkEOb4bed9QWjgT0+dHS0fM75pW3dxjJ5cJ72cyEXrCBD4OBEwjo7h2WKbHfU
2m3rdvRsfqqARepGxr+0QnqcC6yjMGMpBUTsdi3M3Tiu1JU2MKKP9USOtSsC/c1aXdiv34FSdlQt
ioDKYRUbaQFcdF7kewRZmBXIEjtE6WzIuDt2ynUK4gPWQ7n+M46r1GK1WtjcAwjiA0f/rfx7GP06
6xBCxx25Tlok8Mr238pli+vS2elsi8B+U7hJyqkx8iLvtaVipTEdIz/2U/I72XHffZnrkMmCQ7Gr
OOlLvIDg/HjiiU6dIXJU8335aP6MOx/Htie5oQdGl+qm3oopAkl2Mank8df/JKGUiqZ3lBIokgca
UQKoz1+iys/7Zn2/EzYZ++Fzs6csVVR33wwkY+Yld4jlH2UltwOyMcZY3kNxIgYnjl2FCRVGsXH/
jOeiPML/Uxwrpvb4QI9zFTdGg+kIVBmubxHVKZY3F28/yubBzF/jRXiTpLJeYtgmRIrX803v2XZV
VsWF6G9f874oUQl/6IkGSAkjVblFSipqShnSIqZXI2x5svlqdProAMqN2A9eMQ0PsSVuJQWNKSW8
gALovuouSE7dU2Ook13I+pyrbjuDrJwlp67FeearjXVL/m0FAKXLU/F8A0Dn4Et/2dtMArouvrGl
Ytc9UKaTj9nD2gEJt7ggfT7RjIkbzRM12YDqAXOWQMNyeauaxQQNVs9Avq/AL6n6GdAsztWGuFah
uHeSyX6Hj1tx66leuFdqymhrfdjr9EVsA8gg2vLghbvlpd7MCU09cKxghMIke4w2EaY5Oan7QKep
x9UVPE2OcXi6HmtuYAGAxKS7SFMG+yf68oHdLiAs8092ISitTM68yjyt3qxxSF5nqU+uTPtkqXqD
EoHKLNXy7aJFo8W9f/k1InnChlyu7qILLzvuuRNapNoTvpClwoZXcCAGUN8TZyrqnWQHGsVQRkDK
c6z3EC+9oqVrioWXKoZL9zh/j/hrEKcWpAMcNELqjOipKCPKDzGQFsmiVazDO+oDG0ROEkJk1qF6
cskhcN4IFav25YFVEunB3eIJ4gYL77iUJAie/6Dz7IzXlGSBOtwuev2oEiZdG8gT2INi2wPD7Ca6
B8SniuY9+1t5cS/RSYLDPA9i50YjHuW4BSTbeda5oxEsuH7b539BuLUf9W6/UnGj+44TGkHOXzWi
ChPB1YIoyDfCMohZRJsWssD4uSyWZLi4I6rKuZH3c5Y4Q9LeJbLVx5Vg11l0CWffRRcZR1uM4chO
NS9NIcNalpm/KtJDkCR4VpxGtmXneUpBZelPnEHwuG6PsAcmyWntvmxH0g/HoB5l1yNYSSEXY5WQ
wnV86WjBEYn1GQ6Ml/kPZXZT59/RV2W2y4L4rSGTC1j05DSdAHQFUporhb5QCT90ARhhP3ATK6K3
Ckko90olm/Sn+D4En5UUZ6rxDjx2Yw4fnDnx5YMJNQ1Ya6uGNPbsD0ZkSeiqqGZN+2OyBkI6MsAV
RQSZiFAbPS8fV4aB6y3FBZKhz2IjIStNjk5XxTMm7+Ag22HOj0WIpDnuv9cK8qkQ28mgeuqlmqfw
NLPF3AIGkmKtRdi28AN8uKI0vg50zz/gCMcXOPaHlE061z5ypgQhU1hXsH/7Xe0ayfHzLIAizXoV
JLJroqZC8A4iDyJ9r3H1lJg8aP6CSzaAbm93xZ28KInLxC8gJ9p26hVHyPX8SLaS4XSkkCQAZPBa
ZQPx52TDvj3dDHwUphpfyBCloEKL/60xDTts/XoEWKF4RTL5f2P4O7YPJs44AJg/GzYt7HEIjaqi
+Lk+zvg/AWMGvGiWov8F65+DMvz+O13PToaGiHNqJPJV+flqo8t/vCZy0BVToxG0IdFqvzxjsUgH
y9X/DHgu8LzZFr57ElEE0eE3mOrBJfjwXhFEssG/m4O9Xy1w6xaF75IL9eOdPzC9DkF29+J/Svia
knaTUZfxBc6rzB0E2oTXEqEUuc+qa4JmkHWp5sbd7+Cm40XHHKTVj/g1czbzfE5bBrAmYP87/4WE
0k/csIs6Z3MK/2HaIS2KBj7yBCfET/PheaEnDYMlkZgT+c8y1wPDWa+pzoF61b6v9Gun78GwD/oF
B+TIMLAHd7OkQUVDrsrhRVnWs2Ds7DUVtlj6YJbmRE1GkF5apOMAKjcd5uaag3Wqe9aVNxM896I0
Lx8OnsbCMpSmBsi5TdZLCVhjeHE9fKOSl7wKaXpJY6RArzM2S7239Z5Ph1HJ7GPQiBcr4sdRYDxu
WYrMTsvDmXucZJWheD84LyPA83EHONicxKr7R0S3N6GhkyrJDsJcGzXC1nC/bbkExxAqpfl/0oS4
aDODUoGEujPZdwJIitx2O2I72nP4k9Wno2aXWKEJDdW/Ov9cvYP2oLSKhe5f8wh7zawuUONILuop
J8j1zU+fll6Kz/OZc180+M/nXmfhTPhYFI0RsP6AH/XyZPnFAd0PjC+4hrjdqMKMXIgqPuMaz1pq
VO0eIC08+BykIT7+Fz6749W4X0mxAkvJo2g74EuNp31nXAx61CrZ+3XDBSAvoQQDQPfYwhQ7PU+B
C0qSWr8xZfKm24UDvCmH+9ofZOkB4rloe+UWRE6VWBW1ki8F5PsbC9uKSAH8dmrJBtGdS5d+ZcC7
1J3GruY4Ns0yVbsBC7uUIbhGfptEG7P7sXqcacYebnw/9D3yMDoORahDnY0lEwU7D9lOS9mUEkkV
CPyt2duoay4qokJ8zcsFkJoJDwtBoKuj8p0JeJ8U3rMYuq/kmM+7n8wIbCBG9HZiW8QdmZP6ERkq
iduL1MW22/joN+Dmnawi4N5oNQv4YYBTRhgZdMCMIsQh6z4ViYsXE/qvvlfNKRBR3mbwYff+1tgC
xl9ZcQ9veWFn7cbv5IacVOdUX58IS/HXmZwOBLdZuxevz8oi4x2WnzfNAdzCySQElBpVQlMwrw5A
jZ+6hMSYH7xt+Ft+OZhveeBwAc87DH60h7chPuXcQC4ActZVgoXTQGSIx6Gunkj6ILecl5qyEVIY
iKb5GNmUzSxaNNuFpOG/H46P4M4fxiRcXLIi4gR1mvryGHabYBSBsoGVgY58KmSPGRLe2S2pbvBj
9wWy6KWiUE1fqukCkCOMmwBy/is/LcrVlKennaV2qzBo/YqYwxZ2G5h3HusgQuP/hzToK87xXLFV
J9yEYlADtxDME/O/JntY6+vmCYTQRvYH85DxhlQvUNvDSCKg7gFoOTy0ts/RwT/8IumYuEh4/DFI
JyoeAq4aLxVsMFMasl78tbM4/IUspQRzyC57r1G/RWTPr7JHLbA/KEdkjfdUsl57GIV+vKe4yHbD
gsiHc1p0oz+UbwxW942EBWNdq+uGTJKSvkQM3sA2GfqSALfJ1WDtSZ8GiZkI2WEtfkPIEf6xtvjc
6tncBWqChBOhjwlPV03bUZvhYBBZwriOJqePbMG7OmmGJUgL1T+naYaCXVGJ9aTpF6rDVd0f+DSu
EpEYN/BDRmAO9qw2GRE8kQJVqceDZFVbR2EnO53uVdgxZwNskHn06uFOYN3kGc4RwScOmrQkwtEk
4oGVEvmMgUHe+PGUF7TXS/Rq8N/DsGjp83aRUGflrzK/Lt3QT107UoHS0FUGHEavWodpPUlwLO15
vRvVgA4CIpMrhnd+iucHn4iZhGBHO8Avlnk1uXUe7dxfAZ78fw7Rwur+fJfxxAyJwbeo0+cfTfq8
8VK/IoJYoZhFxQ7N2ZAK9zOHDILLE4TOBHLkFEqwWJOEUTdkV13HZdnPF+xRRl2QUXK3RDygYQ/s
gPAYk7X2ccjckR0fflD2NCg/4i+5+7RdavOrqCwzy3vGZLxTLP6TpUqTstaR4NnI2NJjMpPw2hXZ
0Y1sYlAqljD4PRxN8Eb8mgQ4quUGibe2zb/zMN2hA41BfZVglSPEmxwruhzcLzF/6rwKmidh4dCX
CQszqPIHoJ9BHnWai4pFhRnQLG5/ZSDF0QWpQHk8++JR0SaiFoxw35Sa9ENMOY/zXuvDEJCGYAB0
6FmIe+CNRld98kKNNaLxSwG51gV34f4DiRRGKk4nFtgRnsGYoh487v1QN15XhCk427ISNfqV5QtM
FbhpV1gLuT3HoyvuMpA/w7m59pqTPgpRHzoZKlOXi1C45uae+uTuQw4xJyGCSQ++Isg4DV3tLC8O
+4twvx3mUxnh0Yqs8YIn7micvHnPyj3pO87u7wO27vEjOty95fMx2dECoRKn1734UBDFLOE9LqG5
TYNIAIGub/Vyy0HvBOjannPUWtUkXBk23E/IX5y5z7CSVmWyWkij+Exli7cneic+/8WNGGhpNwn5
CRuG+8KMKD770KtetqZII3WLL7rueTL9UV55N/XwthoMooUnfbG/wJxW9YBbyYAHiI6/665kWHHg
g6eQy42mqYgJ8jBX3F8KWR+J72gD/byVxU/WMdSW3fomwdMsZscYTVOtFOjNp9HfpITPODiNyjfe
0rU55RIKM4HrYDLhRwKOv5oYwnRhKTJrKioTso2DSU3NE8JavQPEO8HgfeLx0dE2Ewi6YnNYZ0eL
t4H5PKbbSF6V3SMIoKoxrSFeDZ0/+OlT3B4+mgcbuLl2HkqCF1wznkteuO7pTOvXqQbKTsWor0cK
pd04pHMuE4I3OPR7ABEsDkg089m0seBafrmCnZpsROhT9VBeUVoMeOizbfPuG42tEaJL2qtve4nd
H7cFF/mRdDBxdJPLdaur/+0JWKvK6Tjbj5/1Xj8+Ur6HxgG4L4iiFbK0VW80Hbh18sarI37YXFTv
7G/daZpO50RsGZzgOW1dHDosOAIDtcpTsGjCFpycAm0ePmDpsYYf/b3xW5b5FrePCVpj5PtOcZ0p
/tKM02x6wgla1fYlycQ4IFL6Lao0ixMgW7264vba9eSlGnt+HPi+bhdtIdeEYAROidMow0srJHNm
HuLGNXxkWPZo9iDr/INe13FQ3dFfQtyA9ctQpah5SHRbJZqJ5+SMYM0X2rFAUNzxB2VKprkI3Pua
NyR0akDLEQbhTjgmNlvgkobUN1umwqB/ItDo2+Ut/AG4bk9KoX+A4uxkrVVfJ3eSQC1ld5S8q90c
ErRP0BJprB9fY2Juk5XAztErsXyMWkrXwGChPEIPYbMRdnYVGllqPMW+EJFWFRLkhvcvwHpNUNjs
SYC1BjbrsNPFy2dHuW4hEYEc8pH9W9OOQXDR6Kp3vWH/GkTFw/Edp7dA/5YboS/CDQvyOEQhIyTJ
2RY47Nq8cgEUOk1OAVdhlNOPY1dc4WBWsIbar056Mi29j9QLZq57kt5TB3ih3Jrsq6U47X9H8Urh
Jv28djMdDEe23pRcvGoyafmykFBnNJBjEIgpdKy0OZc+Z9vLhs9mlb22VzTHiZk7tU0DNuoNzaan
vKYPbvEphRBXrEyDwqBL0Rzh1wbpVGMHxBBq/4Iw+ikV7ZMc9kYm6GvHUgpEdpCi38KG0YOlqS2N
QVbajxLpuJfPMAHyE07T6HgU57AveDN8Ftu9gtCWkJBNlfWvieK258P7fbUfliCG2pWw2EHbFzAU
722+AcxEJrFVKDtcDF+zr3Id3v8izb62YYf85lYnBrzaAbTK4snlQ0FtPZBJSF/Vp4Fa4LD3C4FY
5aFpgS3jRSms88J2fZpASxZhdTwaFzLcfyA5pnpYqjdGphHPk0AoZAlpVg/lQOUGQnOK/zBe6vTp
XykSASUUhOsv4W1rJJnb0unOha9PzcVP82/fCIVErt9XgS5MCH7Voo8e5jnSvLbjBQ8eUyb93u6o
NEIzMTiSOPOQ1E5oBLchVnXToTQSsMkbGWIqdV4Miyi+j7CSkxo1WdbUZ6E/1IuNfo+P6RthH8Lv
UaGdOYlu+8x0VfX4hCVTrb/t0ilYOwIVkTy4pxaYwYhU8XxasuI40mvzasnntXKR4ULXj22CPViK
E67kKINPA8N7PnOjRpaQHNm8feFlNJnh/ayV/jYynNvrl/vm2wxWUcqVU1tciQ2rkFPE7i83KJu9
B7u2baQlRQaSDlFfCyZdrEqM+0vH9cfc5X26g1UQZXsSWTyjV8jSYhy9uo2S+BEZSbiC4k5CgMQv
/7/4h/kHGVFfDsP76Cup15z0F2XQPGemEOhuN22gv1jr2UiR1L4uUQ2pJeLdGJyE4OzKgadc2zj3
LxQp92phnqNGHyjWGCA/OYswCDZPHW+DbvjOvICPh/Yw5mPuVCrrdJCMpSJQJziWXs5pyOEcDiyo
ennB4PLjcepcYC27U2SiW2j2pmjNaWpS6Pn1psnMXB4FZ+BLncoUpC57oDuJ1qwasM7sNcX5TgWe
h4Q8wUTju8UQQ2myxoViJMV+jB/5c4DE+L3uwGERyxZNify+jNafc00Kf/dU59mx5V8MUMv5Ni8O
v7mBTpEM/8btIoS+N2CyDZNQxqcfK9wNYl+HSBQACf9SVKNxc+XwvvuPh8WYnMQxPgXuPh9W+DgN
RjMsAU1mqEM97sdpGcFZlaXAen4kQhi2Ey4zhn0svg6cwssGaif8TFikq4orzN3FyeUJNpcd/ewQ
Uq5HdehVOGUy23hsNRvoTIOyTl2bQrnXq0MAZrsoxCMImfY4QZQi/bQfielWXJuUi/aXt8wP1PNd
br8u2e1PKBF6pEqgCUwMuxh6m+mVtxlOCmtZ9rBzFyxnEOWpGYU3DnHaulvbrC1GyBGG+gAosfXk
yUJFFt+jGElUkzZxgQisAyyPff39BGOIIWB8LcDmgYf14Rg5Hsrdcg/OTbdxY9ruSAKFoFeU4SMw
ojY6aZSIqXaiOYtnJ9d+lMkOu5zQQcmtxAgab+31Y/EAcYrIS6QbwS5I2WjLGeHhi1LfmNOg6fiR
qAuJNPw7UHm4yH63Wn7UVsUe7hoOi9ra+p76qJsG2TTuimOouovcYVjtzrlXXeuMqbpLnSUVEcOY
AZOk191GqdE5kGjtjSVCeBRcWoFGHrB86elu0gn8Fn3JpYmrQJkq/TTyI9BURhhc2pajaA2kzv1T
LgQL3hxQGOtqjbB2DGQmMzhkQZjZ7vvFl/wCqLjo50fvSXgUatpdhSa/7EP085I9WQprCpqGyrtJ
sWtikx849mB3HlSUQdrDWV4DbaJJqI8vvoIPmwn+IiNguDMSweg+BfsRGC7DDBrMK54muWq6hMo6
PKPxWJ3LUEE6+D7wNMvTC8LdrUg5WN29ThI6Tfy93311FrYjrmxuY4CO4KvAk/fs7rGc+4wpcPFw
1lWB7dmXHgRL23LrdiMUenp+dmC8XLOXQo+CjGXwkw1FpUEWJkOsFV43+hRlj+ZWsQtdQ/SBVnlL
nY79btNkj3Isv5rSttLRBVLT9vgBOncD13VyPZU+e91+q0Rf1W4ANFFY7iLHpYLb0aSM9/dzoFJ6
vQuSE0mGbxF1RwQJEo2FEfB5dBb5g61OzW2ii5e01a9/FsBH+ehBQjgLPGN8DFNgCVhHZKwU3g59
q/k72diZC8RxnUVT0FBKtWRe2VIQWgtJhWDGEMJPnSjf7rNfTibGMAxbRvlzxyLHbAkrXjUlwAS3
nBzt8SyGNaqGF0tUPwcgsXTHbB4OHGOH9EvVOx5ybyJyT9qpEP9hRY9KdXxAjVicnft2uH9/PFg4
7i5u2a+2+Akn0BnAIwucVRlNHwlFyQSjUBXYAqIMT4kHGZfyJOZ+n1MKWtvXzdccgkb2nPm53+mW
LgLmQ6GmuQV61SLpZsi0JLFWdNtUTHzGB87H+/UfgPusYKXNCeQ1RoNoHyAgPZcbbYT+LKfCwUn3
LPkR3y0DVgMI8B/facJY4EthHb1woaUall+52at1CCtvrUa7AVdk9OCzqYXuv0LJMGIFwDZBZLId
y86aIKuVK0mBmnpl1HQD5tFnOi/nUr5nS9l6GiDCbGjCo+1JNIc4Lj2/OQo65A5UyzveCMLk9IJ/
YDhmShWL6DUIh6j/laMKQHx9Mkv3GlZuvzBqXC9DnTaFs3IWcv9IUI7C4inra+InDPty2+LwGerQ
VFwlHWP7lhrjBpd4gOW9DLZtP5G1hp310KerOBEn7rTSvyslGfAzJOzclt5ZPm1bYSlDjuWKagSs
uIdAasTU1uDrgftRF+XZhS/ze1SITiwW7n8R26LxZHd+Lu5IX4mW6YjsziOfI2Q/VrPhEm4Iu2I4
EZj/P7Ntsln1CKHIepL2uVCi5a+0npC3YeXeepVthqxeTDFrclucG2hLs/4uXvSKu3yrsGUG+ZUL
6FVF5NQ2ZB77QAu/niPkPuNGzCtQ+AJQNGfkY3RT32SqiUX0jUNeFz/bzuW5rtvJFu+9CaJSfZUi
Vn2WgBZ31rMTKdEDLET8L2S6bRK1NUFzSehhZPDD9NxhJ68SbcTiXpqWn942Z+AE6vHKDiKcEOb1
ZpePXPcL60zlVYBmivZ+q8qJLSj46uysUCLXzGZmwMEcXfmxBo4hRH4+H52UaemCAxap9y19YVw5
UMHq9HLeXNrnecpfwXaorJvUemWVmnaC/VZKDEH+yDPLNxtusj8Hcv0N6sZStMMc6plqQDnIaITE
TJMtTZD0L5AmYxJmMjPQZLf3uj6dLhougDI7wjWKybTJFspwLl2/6G515hwHpVXBoMQ7/uDVNPSs
c28WXIIXlNEwsxPGifQO3LN1AmLYEL0cx3eCW7UzTb/K5NvWSIetRnjauHkNxIFFIwT/RUuqtnhV
xp/Gb9e8tDI+1fPECOyc5AB/J2DMP294q4mPC3xJfsZNLlQa27mevaRajTdyEF4ZmhlTspqYmgez
9dNpWAQx5gkCeALBahaUmaY/LW9Dm9owo1j11IuF5JbaFGIXjGRZCafaQTPbJx6zFF+lQ77bE9n0
IK1ZbRebSy/8QGlUJScxo6rpCQ2id/YSC1cniRlN+w2MvJiI7Cut3QtuVvhiPL+57VuVbMQTBfQR
8tAddE/677LuAkXY6AjxU6TKBWsOEFJQF6xmYakh0EC13J8E59IwLFrmVxhLTONcjMXMex/UqO7A
tI7vWOzXGuno0vQRGTLXKQrdn0o89IiSbkwFrHcHROf96aIt8wH2oy56gc7gE/lYvZO+/uBoobJv
+5DBVSeW5TaVBhF1E55481uqhRk+IR7Y3cjMK7KrmXr04xL1NJxE6IvbDE7PJNdzt2xbjXbxVb4O
mYuy+sVWuM2KfWNjGK5t97whl9fEHRIutOS9kXBnJuD9aSHL7hukLJzSr0LWOcsUEPKgmJUc8aR3
ZW0fPLOHF65YPAIYWSH2B21o7a8wWKDy12dKEtIqbI6l61mCUPElrkeUOLnRRbtFtd13upj0ooGw
8646y7L2JP0kA+HfAFVsbAGUvc8oDeCwTju9e0z9LZO7c7LBezimyUQIXMh6QZbMiVhDExAvg0Ag
554NkP/kzwwDBhRzr2D5J8OEHUWbkjZA9dGB/I/mNBJ3plswUPZ8DEJmHW5rNmT9UE8X+h9hQDkS
gED34cyxthoJZesqps8bCRtdQ/r9DY/IbdDX5sdyyXHYQhRJyVt0Nj2euwYsv+vvpor438AIC6gY
M3xnjgk2OxwpXDnJqOEJjIBdQ96YRLJblvfUQISQ3Se6GqYkcJqurEvt6Hns60lgpjuRQMlueP2f
IPZ05OJCfn+BbJkjGLkgd2pFk7nfQ14/wSyaGuwm6B8r9Ld1BprcVEYxjsygUy5eCWloXOoIEFJ9
jtKmEZOdNwHqM/tNklgCX3xs6g4ScVtl/tATb8jeXtyrI7v3G5TXdE70olP+lV9HLfnb6mNsuWIM
KGDKSRwxCzNmsDCXTUcyD+6UsHuqRCNZ5fxiDcQUiznIgFOLHJXRTk1mxhWCr/IL7hPEpcI9CK+Y
ajmj+Ly9T+RGxyjDpGumrUJqkrhfs516Yjq73w65f4xesCgZfohwNZ7JHE1yEHH3x5kcyENj5FFs
Nla6pX1K3JahXQgt0J2Xl1Q+Vk9IuImmwBbYTmVMFGc1ScG6wZ/ag3pm6gGkQEPYizyvLYZI26Rb
Cfr/PX3zwW5aE+VAwCEdLl6uBACe9I2MKD4lS8LzmVCuSTtefbI+8LFFAhpHGd9/E5niUSGWHl6g
QXNSMD4q7GGJ43Af/q7E5ujA8zMJ8k2qwQfrng+MQfC7QR//QyVlhzu33C7lE25h+qIIAeo28/Pq
G5crV+CY+HaezgSynrmSNZWfuUXScEEiknAs3Hkhpsvw7Y7gv89gDMRNX38ozgNjIcIdCN0CbH+l
8LjZ/M0NNZ5jgwVWggvA3LgVq1QxU8wxoRE401GiOB2SV8ywVoUhR1TLnqeqIHQc3RwPAXpBGhqd
H1txW6u43oYcEwlfnRUblDShsok5jJu1Gl8vWtBRKfG7OhWRcwCjeaBhmX++sXpVWdPhdXX6wpOH
n0GEv0HDnvy9CuB18ahLD2UKvCLb3P8tFBwax/1kKbK6ytvR4z2tOEcirMJd5ajCChpG/LwxTMXM
BM5GBlO/uzpWPFxmbDOp7Sa8InTFHVAAU03W52rdqJCNipikYxJ7JLkuuVK626JnH0lTjdQ2yu0t
vFpx6LdShvxgcxb7gJW+vokkUTAr2iKG9LWCziZL1voCO01PRlEMPEWj4njNJwI0vHojhRNbgGkl
4TeQYmx94nn7j8k1hxEyN1Li+30YZV+/8CbCL1WYm+peEJQodLzED0bD4b5+8ZIpIXTjSvHveEx6
zZhBpYNxaiu4/39eGoPPRyTnmLlLU5GIb615UhQpwdxIPcEkVFP1ovlMX9ULw0oCHpIW1cL7ow0v
7VHdeh623Lkjdl/BqGnNNYbEDTpRJdGK6432MolQ0sycSX2Xmd6KOyA7BGc49Jl/m+MKWQOor2VB
RvAdAU6n4C3/SwcD5EM8msfMe6P0prxRRX0iYiGLBKu0GofZeb4Q2VY+dQpBzjVObtwdDe+ah5ZV
KYEsqQOWGbjYcUhDjdaC7wTkwEhVn7wHDFSSLWtR20MyCeGaXeVAM7epchAbndpgwgR7+tWPOzRf
FIBLD6I+TLc9mZveFj5jQIo/qGX7X6+jb5SJZD3p0ak4JgAq2ZGf/sYJZx/kLlm4GcdjO1U8Ur6z
BbFYIXczsFOCgngBlIo15iR3zyogjk5t6tJtOBRQpAWN/ttdz8vmzsdRJ3mjSckDP+kEnD2a/rNk
PuMniBYgIc/REWpf5gCOawTEDT59HsPbx0a2rLXk6/GOo/54cGSW4YZvhfi70sakT1dxDMMNKyDp
noIB3GPGGspHnpKOTN80oJ1VG1CIIRQhsDKVZxF5F63IrEQroynMrP/K5Mea3qfpEEVt9TK2azJc
R3ybG68CbiMKXGeJWeJT9ezfPZy8ATA+6c3v+C/MmRogzDSH8BN3ghDW/NSf/+reZ2GgKUfYK8gI
m1UrtWX0/MsC6WHy7tSa0FWRi0Chast3Gx+eUUzyLYyY/JbC0vze0nKObx/u6X2Kp1MP+IU7/71q
vlAr24XgB+xLP9FFRF+ElVPyG3pfO7hjqqW/8InTbKiGrmch6461K+bDsLZ8FftgsxIPYxP4UT+O
d2i2vaCO2WB0fc+Fg2as16qA+cyn2kNPPt1DI0qAN4S5bZ9ksSf1c16tFXdPE/7oGUFvJX9tpAOd
BG8Jfon1E+4NFzKfz5a73+wrkZwU7ldadKXzPIA14ANVxraDSu1WZ8O7K9XrdluBuV+/CgFmpVdF
QJD9f9vdejYj3glkGDH5lsPdthBUnlsJdL+TGdao6pkY/Gk4Qh+RLtbF7WJAwIf9p2rRXkImWNPi
xRZ9ArfHLWWNyJiqAIvCWcDU8n6qyPIsLU1NHE9w/mPnQuJ+1CQ9K/+QNIrqoeVZJb5Vsu3leW62
KKBy4IaLogbNfx5Y1Vo7q50YxoKzxcbW66dAmQa4lAIi+yxKb+Et+RU82pwZNQq9z5GfKA7GaK4/
PyqfcMjwuMqPpVvq6SARF4XQk16R4IRWyREpTdA3/uDkfgzm49bo8D9PaqHhI5hebOH35eyS/OgH
k+GjnYUmIJDYPHers/nclwRbAzjsOsJ9XMNVieSWSPH+SaisZo1LtSupdRpxhSu2kUqhxdcBgKxx
5MvgLeI7zWVmEnY2EK1sCSjNJNQpQuRQfYvFkbWLeSrZwrdB9N0e+6eMWWmWavjlAa4AX8oeRRrP
icKne7MSXHoDGzqXHY86SRogCFVjObOzyjXJQnS5/nCrloD9YT63iyiWT8e90dAJt0JGJj4lgGGT
WsX7QgSdcy/f02SIZWefkpO8AZQCIGXHzv/mLZUEY01ykYCwZc7Y2S4OhkLTdB5KPCAR82QQBhOD
u3SYN9Yc4WBAO27L0exKVknGT2ovELM0PVw7xMp5pizNB2qNBj96vHUbPsS5PKcyPg6tQMRThPdn
ei0dWL8nGb9+bRdhNozvxvidW6ZlMj2atCX6lV4JBo717J8fnzRs6XSBaGEImtonKqey7+K55Ax8
TdxxTT6Ad8SlP8eBT8hmslSqqEvy4x9itaZi/wqXfNQi1dx08vN6AY8chs3pyLKfnJWzCvpSpiDc
5ZVk00Um+ZS2+nSOYywEnXHT+S3BJWvHe13AIjzolU3m4ebo1jExEGHPym9NY69GdWrGFZBTlMuv
BGW80y5Ik9v1UT5R2F86+Kur7L4trya8cxELNb9ouwPmTtUy8al3Dm1sluXgc92LIEyM24peSBpt
TeVtMyRitRx2GsaYaww42GMtMu7BaUfeVabrrKzRxNkOtsx6c0K+8fmay+TlLjCuSjUQBN6roW18
sF1YzDj+dWBBQNFZ7h2/o4M0ca+VEJ9OauL/IgQsn2bAUWwnPVYjVWX8tDmr4HKMp2IqMKwR8Bhx
5XnL24DnkO6YT/Szt7fPc9DSrmVmEk+ZZ99ujA2VgfVkJSfbsBkJuEsP/vRUCeEVgmV6dz6+3fWK
7WnnYvrEsJo2RwtWKE58DpwQL+5NjNkW+VKE18yXU+ott+S6nsWgMhjnf9e3EkjE5uC/NDlS4axF
32RW3fC6n+sM2CSNLBjEpdSaZoe2saL29l4MJBtVHGZrxy5YHtJdggJjT7Wsqn0HC7Cwqs+FIMJ9
N63WkJuMqnxGarJYtXF/M+sP7IFVdlVRK1hm2PFVtYQVLZK55FmCOZNKWCoY9JeIkvuRE+Afc9PZ
usQE3Jc3S/nK5MrcUlh4AIxTr+YWlmNazWs9kGzJCAEmkAcVQKi3+gqiAELvdYhX+GUzE7KBbH9t
5XeZZIGv6imnql2t62dEx6sXhRpzXPIcjVMcOJI5vTr3IE/6XZDOFcUWhUdiVlLqERoONX8TKMvH
C5oBL/y9nuC0ri23PBbZP6mQ8lqvTUv7Pvrhh6S9GF38l6AtyypWAsQ8QEAjdOhN/QNHV92eGDXA
h4fp7pIA3twzDvG7w3eFOoiKwY9sb4qzMDAbn6Dhx1H01yxJg8JRGZtZzpNu632yM4hJs35CsNou
qu2ozBBbS6TnikxYERdcWmfKhtQ5GqbH2U9YkOzuKvHMvP5i7Gu6KEiL6u/dhumacl8pvHC9aWTH
PfqI3oba/5rbWdWHKAv3571QyeshhEOMMZ1P61y2/75hrRnLRzVCLcdFi/PJw3dImz8gl/wRJk7L
r/2mKdJtez8TDZx6vCtRcLP/tJvMTFbeWq/zehiYRYihsn4CKjyO1WawSO7SQaO/D+ZHxMiHhv+W
Qc9dlVlBtBRokIPkjV+0a/246MMSVdsGNFLiZHGZontedBw+65hZE9xOJwij2Gp2dFkvQ4T4OMQc
rB9K/aGkKArGVBzzBy0YBWuIebHmJbYLavhsUtXwc4cQxKSJuBYXhlruJXZtjW8vSujdWiIQfbp9
A4wVgBMhjQEUtpOz4CugLyN3eNA7/OuJisTFREn4HSask4y+oB0W9wYx7KoNBP4rGXAbdssRCAgo
9VC5ZqCexbC2fdkChXwH0vtfiLX49Z5bqW4InQErmDGbbunyN1Z++Rs9jkfXpHYApJZ8udiLpSOz
Zf5wkQPN2f2hRONXgBOGS73Ib9FngLoJQvQ6cyk61QD6RzVTZiOwI0pc2caKKYOcKVtqG0ktkPBb
Yr6MkaaBYILAznAGiA3itvAxVdb7/OLexkf8daYMFhDXA0jDZA2DL84iVuk5goJS1ZxdXV7+FI7a
/hMP8tIxYRPLroMqUXPvaJDakhukVtPUZJ5j89cNFcf67wIQcTDfmnSgPmbQK/RkVYGIkp/bvpm5
fiSsAJD72M/nQjLAvxUDn+VUjMhrmeeK4M390kPEdqvDd1+TW//oKQTCrV5gxMU8U/V3sT1tN1D9
qiwoA8VhzUAH4Pxf7wm5yVOqkoD7d9wL+mYf2nQ0sQ7JCbDJKWnYrXNbzP/cGSymI1qJgvyRVPIj
fsAJLJk0SQxZb77XyiFOp6h2IwGpiMQuWuXqxO279BeXt3k+nnlnhma5AiAWqCWHfbLzYtwNjyhB
m+WZoLe9XGIFbH3XHTri9Q59UMn3bBvldwz30JgPG3bfL3ziln4COGw2gqUkASchvFC/sX6tUaQD
q1R01jF2+avSjB8XogheU92o9MSYTfd0DM2oWPx9oNY1ikZz0HrBtnH/seloRkqlRDzCB1GoCP40
wJzRYrpG0TE7KwEBD/nJIKf7j2OM4BH3683caLKA8FjbyzaCGkjcdy9RoU3v/C6TMwdsKnIClmpN
725tFiyIrDnxNbo/cMTkjM0iTI8LkD3prj7xHRv5ch4j6l4vCndWo1mRCP8cnHdhzzj5g3oTEnvA
qVUN58WsV1h/K+CO5Rz9j4sCdO2GTk5Ie0vZQeGfX722iwsokYVF4O5M0Ms5FFqo370+PML0k5Hh
G/y4fEEYy/5lBrOT+Dw6oRyFTfGCTMfLS0b7iCZ5rfkfY8IACr8GZivEgQBWuabsz0VbsWoYqu2b
ki+iNv4ExygWSeQ0H4l3MmvMpYXY8X6Rxlv81HUD6uU3MbJ/CW9RUdq8JUeAr9c9V1SXoSSqpSKx
nTfltJncS8McWCwRdOW14Ku0gbOD4IIN8uU0Qa/V3wCvJ4VMudeddHjbsbd4+ayFvO4o1Zu+/U3p
4CS5t4CMroF4Pt5rUeT8hKd/3FaLHXaS2WBYBxt0Mqgn1YOSDin1ENgHF1ntYbTfFWLuqWa52JQg
64zDEEqwAMt5Rg/1WQbDIBe8VgbQ677lpGK3n3zGGh+o75iqvjeA3tjVXdABievL7L6K+CNFEe5z
eohpm/VXh8SJv/O4wWjydGY7h8uEyOTSBfC2P+VBEAnrg+eJWUavFazg+ET+P17kBD16GrKfajoo
ew/TqW1p1YAxQveTxfcQrz6L1CbTmyGmbtL1MauOFD/Ucc2qqtVxjp8NtVg8bSss/Z8OJY8iBSYJ
s3WU15cdIosOAEUKlSDJmCuf2aykuUn9LnkMk8l5OFxuGeuwm99SNeMQOFhw9PHHQ2rZdtfduC4h
wBJARm7b7Uf0NYXAG1MGXGkeeqY3hl+3kP34FAAdH2+/4KMfEvJIElEzqKgjOG0WYbYwqVZ7sYKe
FmwkBsJbhALgnJx0+bq7P2JPRjwqxN1MdAliSE71IxLLi+5w87xo99i8kZJKBAP45bbBt8qYm13K
kzk6fmSNzYdvIDW9MXMFTxUCITCbjb9Oa684+GnKY1mPlLUYCy4n8YxsIebwBIKmz/CQCtr2BM/B
nAJBjCTML+uEjjf+VH7RSVSsJioXQ0AZsg1OOD5M9j0cFngBQOdgf5coYoENsp1YsMjlDzn8Pir1
OC/Jbk/y1Mr87MDjHFyFHdkkwZBFFAxjBnQMdOtcw+lN2SN0B5OP17OgbsPOPg1fFgaPgfnPETjo
o/iDyBOhPrnvgKrI4Ha63vgwa1TN52xQU7Q+jCYlVI9QkqxInzuITLL5KucaomQkaGcQWlkY2NVB
lJowaaVeVrw84x6TpVY5fTK2b+cKcbRt/qyIUYt90mKGIONrTwzstLjQDYeHQu5w5WZGydeyTGb3
D16cE7XAyg/Tg9G1fZqUctvGHDK/e1BvTapianw4w90MCzr1PZmqzNBjjhUVwRWni9BsGG/nptaf
lv404BBzhEL6j0URTzME7WF1sWUvB8vcEAEInHV6pjgxUI7hR71SHWZ/prgycng6RKoJUjciPOkG
N8g/YejqjipNRUCaToEIBW+M21dMu8z1sX+Gd1bJni99FuVOLOAXjFbUKLRsZiGWah0QpTQzvIW7
z8g2bJqp8QSkNydsCYGSSdk8xYGsYiqR7phmC7gZeKzEuwl/9xPnixnmjLX0e3sca3WwcHMU1RpN
T/1nchGThS8y7i3lnCA+YhiDY8xN2pJjOB3+8Tgg4FpuYjkHOaKBGO6dEhfjmeQSpNL0A+HWvp2+
5uazQ7P7/P9hp8Q882jZ415SuuQs2B1hzmiT8aTBxZlFA74CyCwwoApr9mBAGhxa/GMyp7P2F84j
QdM6No0Wv1vFHIYthSs8HVNI50ZAoOrjYBW/k/pIncuvEimHubLbDxvVPojq+mMDm09e99NXA0DN
1uU16G4LyPQ2S4WO8YLipQRDY+W/n5ibSm2cYFQnOgSATdXNlblJMhZIiwS+Yg9y9Q3CPUSpXvdx
RdFwm7PNQ+WLlMYkn9OQXshpI9Gq+5fQiqQlUHub1PHJMLIQknPU2pHPQdbpdYk/4WYSMnSK/uMS
PS3fuefN/Wag067OvJlYAkWu+g0lMR50TAD18ljhDvFoKv5k6CHC5lhqlgOZdCfGSPAtVQ0Ol3gj
G8NI6J+yj9YcV+VEyyEvh6+yW/pDpO+64ehRboUH0L3SzzvEqD1vr2793zZoaT7LWA2+WC4yY3m3
TMzzwUe5tZQecPW5zlZFs0OL02qPvrvLZwy0yawiL5RpknI5L0xcPcT9cIDGVbpG0Sr4/N6qfIRd
gmOJiErVwi/xQ+FOUlAJAq5lkZKCGwlzB62gCjVqsoK3dvfk3bJpa084Lplq5YZVQnLNcQCFhvP+
mgh871+/Xwa303LmwF7Y92C4xBA2f4L2+Xty+/9lt/KF3SAA2trg2IrIAmybjbqf0557etz69rQC
4z0DtOH4nGFZGhealBZ7RIP720mpvqEYCx4t2me0ER3m6LAAEmqVst0WIAsY5kdriSyRCU9rmOpM
WmD+JqGIPCzqzDj8id5eQmBIcyFRBf8bEuBfAtla10yAfPWERKQvb6ARAhhoAvGRtw6iPvpq7VYq
GZkjmkE7nyBORCentGQUvkCr2KzC8+kh4R4zLlyVK/fOZ0aBs2F+JRIXWDlrl1Wb6gUhnZiBY+W9
WBBMzeVXJ+KzK7Pq5YBzqFaEj8BN/xdM/9UGQ4Thi7gEzguuBkJpyfR91t38NoSh2x5rHCeMio25
TfdkK2cyVYPhPPkmhQxY5hr4QJdXeME0NL4vRXP/uVnVaXKMIUtgUvLP9aiFDSoHVmnZF0u/g92l
nW/EyHO7HwvmDnSOjmu6TAsfrzu1xvU8fx8d1FTbSdI0WZMErkzgUU0n8+FSQU+vGP7ttYH4tU4L
qm0+d9TeETtMnmSF89hUPPMRwX6WBsWCiTxq2B0jnSg6lG6JCIlhPltCNkRcyArfk0ckU/R6xZZ0
xxVBtk7bO47czXCp39Q1+3xOMBy6f9vI58SgHUVF3qH2RY7jlrNayX5v0CkVfCkovlBuVgCADfRI
c6ykUhwBPpdScgFWXSzgyH+Z0gHHzl0IAUihmuwmiduJl55qpSCSX+bzv+0jhFk3JLECgjKzAJMw
g5K8PmTWx5lFy6j2tKVUaSB/oP5eYDkZfxkoua88pJZCHk+kbTTLL+RgNp3LneQOhhkUlakXjAKm
6dpETpBX94HaJDT5eh7S1itTx92V+479S+D5/7j9HUpRzc4xep3YWc4jmvNh3zLQJsTcWdP6r+LF
e18cb8lBtR6/FnAE0qQf8wULO7dwAm5Y5AFvak/glCUgtQePoV+wHBK+qmOS275NVYnvUMDYnzYl
ucXCmzveg6J+FUQDG8iC7Pl166O8IYRIFQqxNoBQUgGFDIZg+xM9yz2GfuiK/XLTwJ+gUp/0rfuX
KeiUDvlhm9xeX2mlD71pnwdQdnFktijF2WY2kuVcLsgA3dH+UDMLg3QKE9Ni9EVN/ErbASuu7O/y
C8njYvuQ9rRiADIjP7DXsGWko++m8nRsVUu7xdVs67DwIaJ3p2DrzNCL0jpHb3+wXNX0IaBSTsu+
w+qAPmAP4XgHg5PZwlQRMyPw0+y5fq108gTqhsJfKfsxaCsxN7ijtt9KWkV57iwb4CKb5dr88WSD
/hHh+fgb/K1Ka7zUH9ohE6Oedal343+sIGQmqxa6OqkvkrdMRwCEDU0+bZZBwxobWGXrSyS2cTa+
hyLmeX7gyqla+Bpf7DORz7NAIKGwkG3TkPCnkSfqHrMWl7fj4eIRx8Pbj2zd/zCLBoTkjRhHPFAy
wKTXBqbYaWGYI9DCsQ8D/RhAOTsKEs5i8XKsd7a5wwqZmXbLLQJO3JlsB4GtvRyZVMmfGuhPozD/
43C73mdeJDm+ePkakDErUENvpMDPyH6aoQbZvwG1mr4UCyD67WgDqqj3z5aWYpxS2643ds31BoY6
CX+0IRAYUkXq5G1qExz0BQk3FxJfunP4hGqUt6TxEHysN26j7Nc1GyGg+Rs6htkjZb64UsTjKYI4
qvs3NuwyL3+a4Rvg651lOv/ZQGEL+fHu1p9HSJbk8z+a9ghG8LySIgJ3GJRQTivaeoW3bVL3sTi2
5I9h5e1i0eKtyGzk3ymcK2gJRGXinj1pfY111KO/DW481qZwyf8sidnKxB0VM3xIRmwS57wHSQq2
M8V6hpV+XY8MFBk/JvilxuVR204Caz2ajsDpaMuIoT9tUrkzj5UQ7bDIlufEWTuuFkLVG5GwfzgM
ZL2Y96+SydvtryO7ejJMtL8wLNuf/rirq/93FKe/TZ9SAsUgDimkHtEN2e5wgoFsWPGgyac5Sn/H
iCtllJFZVirbITiDuq6nFOiTXhx53e0JhVv2nmyJhcRxED5U9vOsURODunJO3jCNVdxcK6tSjuoA
QML6AIEuUkL4+tATwpH/pPxt0wt1gkO0M+5wa1lBbGJQInCwtzMYeIa+FQ6+xldjNF86DRt8iz92
X2x4Qz1ziEG1aLj0AXoDjwKFBL3NNFUdoYty3TPG0pFDuL86sBYPQw2OD7p5cvJla9GRfOdbABvD
DHGZBTGbilkAi1h94MecNMB8/yqJP6L3uSPN2UKfgvjPAGEz+AGr62hlIXY2E9A4UK+0pOlR3num
TZGyoeBKGGD69lsWti31JYIDxubVxqyQVcFJ/QICCz9W0kjAmPCDXGoOcbdj8vTA0moX932KTatU
yYdg+eY/WoBwK196pAzU/A2qN0zCJTfrqWztm4tkT7g/d08B61SAIq+MoR1KacwjrgDVJTiuPSNd
Nym+D7937s+/VvNGmeB12yvJeVF5q5j2H8OZQ3MOM5mnL3oS+2w7kOBTlal3+6aez18eZbCBl8V+
HUUsL+RAr4yff1RDLedNffL9wErG1//FSMyk+r7pqqzuPrdZpMddGK/Vq95WY/5+s0hPqpqrI+gP
LeKLnfZX2WBEC7V0vLGI3WypI9h5l7j6kYKfDPpOBonAmPHEIRUxh+xYGLglAV1ImdxLsm+l/GQs
TU8HXlWEU0FL6RWMZ81GrkQ4hfRPifZNCaeN79oYYJ7PDowhhipleDLmfOGjKQU6Lo6G0gh/Q2r6
rD/c5WbNPV0xNHWr4jSFqKhMD18xXojA1LhxRHXdbibvJEqvCLyTnOTW67kEeevr++xgOnyzAPO5
lpiocLOZrWhgdwFyUVfxGRyXHTwskSov4V3lPboOnQby9+R7yig4OHXX/tf/xUcAqOe53Vz+mmU0
9kjuyYfJfXYEDG33RPO27+0ygJTTlBvcFoVsLjM3zEBxUeUuOgWXz/CKDnamd6qgEi7x3vKodLdB
1f4A9bDCxSTbYuFqn1thPwAArB2QmDCMJWoIsqLhee/Zk3XLLabidd2ypPPj2RfsZUfX5ZJgoDOu
GNA5L8UYAvDa1OHUld+Ue37Pvd6NP5vP72BwhRZX16vothpVGwrZ/HGDgaUYm8r7UYVO7SDKn2bD
VBI9WNjI7QI1uJdGQe3gW7De5TUkA7u5IGkHj1q3vnOwYzc2ZKNfN+2HxOTXBxyXqSuhDRVSHhLV
V3tEDuNHb/JaJ24AzUo/rnhoccDt3IBPQAK9TShipwY228MV5eqfqp0QTV3pYM1tA9aCaCFvK1aW
J85HcjWcDvK0pCxEO31xYQN1HzJzHoAuNtDdn+1Z+0my3KZfspEPyP0zzPBHgVeu4lnsAMQZ6M0J
U31nB8aABLx2XtavCiNEDmqTQZ1ORx4MKnBPhJKF3LKjbd9AwDZRAqsZGblc/DHpsXNrn5cp/t46
rVKrjjGSAXYChuPdA/aKZKekJHL8zRRGVdcxECJQJVN0Yyxjysretm2W7yIu4qvA3dWCQGdfiGbE
oxxju67AyUFzc1zCVIFLj4HIKgrMDWBB1Mu4G63J+RCIb4+v9Wm3/d7wB1MgIwUDezpvmFB1b+s7
LfKcmN4VLDnMvQ8h7Nt84dviP7IMwsYuHTWLMnGir7jqHwKT1hvONWqAAZgQQeNENWCk8sJuYx9C
uqEV1ryTERiX4jC90LlQjN2b2x6kgL/5n/q4EBG+/52Q4z8yxOILe05XST+bpRU8vlXOJbdx7xYi
lGd3nIkZHcjVCFzFEke6kYnftOEV9cLQNt4limMGdFpBOGtzuEOKt88/8pdP+MnEbA3WXNO0vkuk
ByQLoiRz0agpP0T7ndQ/ebP/Ca1KUfeIm28R5r1gyICn0UbK0A3qQiivDoJTuOa6kYOLIeM0rkFO
CgiUWihkG87Bz0pqte+6rFBKvXySj2se9pJKRKdQshjKi4XoW5g/4Y/vP2gO6lDaNlSUL57Unr/W
LAOfbN9n/e5OrNeVIMPxbQ/yRfDJdiWyU2xBVt5xq/64Kdqy3cqPg76gtGsNCWKIznf7BZ3e7BVf
pElbCTNwErpdhnZ9d16ky0eoIU8E4e37vIotflQqeO+EqyPol11PK8zdtJ1uwBt3f0/EEmLxzOlp
Wi3cYN5knu1WALAPE/y0QF0+tO/1VVo5xe4j4BYIAqxcJqXGkHVvWjnoKQ3JH3UmfYdn3cqPPrG1
18i3ey+8viadTMxJ8YFyPbQr0RTNak6NO0h7o2Rf0A3FLpOiw1eeHSKaoKip6QPjEoKvVNtaDWuM
Cn/JD6w+0ufEc2jwCyiyJJ7d9x1P2c4YGXzAjKqvqPXybXoR5PBZc6ssOUfRx6KrSQMUjf/wJmKH
iJS2P+jN2kBTRn7fEJbHKh7SrSRpmvZ2iNNOlhUlzcWqP5dV9aFzW7dt6xfwMVMEjgIm03Q9Z+Zu
ik5/mIGZsxcfl+rUYtMZYmsvgZvjw2U4myV7Sum1SP8PTqT1K8wfte3Vj4iOajaqXsz+QsTNccsV
tWQHngMmxCQVKGFxzawZ7g6psyUoAaJl5oTxUGp/8XH3s5Z5rKBDjr6jU7I+OclO+hhX4R0ggeK5
DUPfXZqv8xlvFhk/yrvaHP8x4ob69DtJl4bSgBn4hb+907SCD4hgcDeug6bT7SoZfKYhYtURF8bm
+cfZoxy+q/4LtT86YWFCwoXzPRmT6wrd26Li75raab/cZMAaEHLyXZhxFvxxuS5Bv7l0wVOa3F0C
iIRgtLkU4QaD4EkkBckoYVJS7QE2hIHOTFjgY02EdSKB/Hdox295te9r8dbRDQBZQ5Y6yR8QXGBY
YXrEVXx6Xaw/52pn3nVqBa/2jipn23ogZHsIG65cIfJi8Ssw6YwqcWHN9EzfIz83AN/OxC60xf8y
mEZj9+pQspzsXelahCdu3qgFYQDKI5EPxEc1EbN4kLsOasucIwLx+LB/zIMe5QrAbDwANBS95lun
xMpxPmGKxZLEkAC8b/XmgpbJDi2c+Mf2set7KtbKPp/dQFt0dGM+JD2KFiGN81uwnxHhs2QQAyrm
7F5cynThAh8sTTg4KwCSPFVORe06mkbeX67jkxl/EBEGeU2bWDXiAs7lbT5C67qhb7caPlevjAuM
JIW9nEwIpO6oQ5uoYJIA95d1bSmj7RfpJ63s/UqYaw5pv01JsZAUxPxiJ+Xj3U15CQUz2cxS3Ggg
zejHvHhUf+WUs6doX8qRII6oj6kASvaA2zQEatz443WxEeb4RWvOlnux2is2P4InZiYppK6WooWM
AH4vkDLHFhR1Q1HrzhOPlND4yADP9qwd1naNDCW9ovksjcnQMCYDQnOaabY7eb8H2MSXcuCgqptk
/618+sOG5k1CMnNGFV6aLTXyAl3KCBb8zoxyxpnlWSiWRDDBFagazx05TAy7JdHOnbhAK1Ka9KsB
QLNObiS92BAUFB9hy7GKyPtUt6cOTXLSfP6+TNBbETxYG1Zhj8q+AnEJLOG8Utpz5ibUbV2SsBSX
5rk7OCH/i5a1ZB+b3ItrKK1qZR/tFgvCXWWA3QG/G+Qz3Jfv1oktKu8BzJU0JcdAZInFElnlpOvb
9LiMPFNDcTFH6FMdWdp/GNgWHBeVAfUJ5Gh+6ImK8NwiCmbrmkYXrVvQTXjIupC7Xl8fI76Q1GYy
K1szNBeQvgAWnY/8SHYZbEHIuoB2SN7KaPQOYTRPUFJgr+8371w29l2SiLetU+X1kJ5ptw+vmJFV
6JZbu18dXtKargY8JzWLN120EgmxbxcQ4olkWdotJ9wA04yUhN/auRdiYTjQDfHMeocgFRViJXo9
tCdEmsTxTUZHpVYtXBwIGbvfSiYEJA9SpyFlsmVlDZdh4ErxsJFmpjF7LrEKKdv5ecH3meC9fMVh
Zq3uvY7IeP+f9e8kUN/Z3f2m1kgR1FegnrNdfrlVPy4Qkx3KAJcha8edGEH7GOqXyUqZXqRK/nSk
S/QcXmuxuD7W0On7wBSqV5qXuN0f/XYQU8alKh7T8XhCOe1fMCzweYn+sknFBdThasNWPifyGs+C
se6VLq8gKo0/Xxzvlv/mqkCG4bHVjfPMo2z8vayy5sADUV14DtHl1dfx7qDf2slNrQu1Dzj5tWcn
Ik6G1PoUTh8NWlED3dGUQ7bZTO7i8y1OwiqVAhHg+dpuNXzwKLIEPuCLHZQG8PZlnbvR2g5Nz65r
rXmth/iyQ9/JvM08iTbpriFJlyUR3cdZFYtcyr4yQKqCRyCbdfItReyEBdi9Y0ZUSScCTTQmk6cx
TTPzomjmA31o7KhejqBk0CSjxKtJyWXDu1YVtia4qVR5HnPfuDEavQhGtyEw6zP/8pRT27jfsvLh
kGi2qphL6VRC/Dse//xU1W5+Bi5QsAZ5edyIAQaOBTzoe8Zy0X8WyXDVK8O2WYWAYvCwHo97RHs2
NQlG6rTsssdesSU7T/lR9Cbm9rR/I7Dez+sJiV4BQO39D1U/trYBl5aipUWNsvx11/O2oyDQT7KE
vcGBsXOhQRaUZ5oZ+xpjr+IYZAkodO+HG5KqNXo3e2n3DQotTIi3JI9ZbAbnOEyT+/3a3B1bRxsE
qlWJqmwLL3bMfR3YB69tKeAmpqtFwnIvpDezHcwUXspjrYQwcY7z2xATMl7Xi1o02AYl4uo0RVsl
EZf95zzpES4CmTUlUeg4VqkWdtsjaZoSBG2d1L48+/eNPjfWAlLHWR7RPiESIxNb6687YXMVfXSl
OIqt+SPNGIviIYv/txiXocEXDJcHKc/SCE96zZxoSvNMtn4dtmUd8vcQqXCsfxfDtJdu0N5VCJni
I6tWa1RMPKRGC/4rsM2O0sMA6P0jEkSMVOG5fiVkss20xo//eIZRoYXWoDhNUT1g6WsVldqXyZ2v
dhjZUjsFjFZ2BNvsVYe5HUA0mmQYsnxw7yE6XAnzcKtP68kND4if+N6Yc30Nq4uNlsf5cBDmiKN/
lY4EBhNDE4M45ZFLmwgIc2gpWAOj6G+xInOONwD43TbGWWGAI1p+4vGNAY8LIQEGkYOlF9T87/Po
eWkY4DrdSGRySIbl0XP/kKQSuF/J8rscHzrxEoouPkrQPLuSjdEsx/CtAGNZhNSGLwn2/+Q2Ye1V
DXjWdBCEGdp3kUlIfcoE3M9GE7+SO/Ye6M6J+JaluhPY5SDKvatDB6LQVtN/uTRHy3oEZLY+8g/j
jERMHlIcOQdhp2QRoaCRCQtDAjK0PRB8whXoGKsnje5AvCkbsEJdXxNqAnJu47DTx3zu1ZjYAJd+
nZqdcBe3R83baF65gHScBCS0HPocM4slVKi8yP/jnuZX5fJ4f83MbLz7GjL2WBcubqZjfgnuyqZB
hlWz/iKYzXrziA8KJOJFuablb7nm0g/j/CMEgSBhU2DnKbUsx0lUJbTD6w/pRl/57mEE0/bRzt7r
UzLPnzZoqlVREuqh7zcKG6WEsnefkHKzz+WjJaMaYfyw0fxggWXJyctN1bhUu+62jFCnABk3ATxE
ZmL87uzPoDyD4B8W7EKLh0lGZF5UBWMtJ6/WyxW+JZyLJRRKN72Z8qgd2dzv5eEP/cITNZdi1cCC
FO4W7fEkBTvxN1CE8vp12ktMN5q61cQXDv5vgiXgJ/MUcNRw+5FEEqhMf179paz387QkBfaBbEaM
mmulmawA25l0DS4JmcUcmAchkyok3XIRsOyZ7BpYrSdOV+i5iXYAHSUZX3YdS44NC/3JUwdCgG+x
pEQGfP3PA0WucuAf5tuYKHUUZMkVLNYSBM70H8AGtvkNVqVieuuL7txO1bq8wWtr7+N8UyKEy3s1
kEx9zSGG6d+MDyabKtRsSUSt8XPAM4lBp4l/je1wGCOCQOTLAWGxQ6HapAuiJEkkANs9Yde1m8lu
0Aru4wS+UvFX9PikSbltJLwBIkHys2fcwNkAzvMKnyvSyS/YrJQ0DFY4tX8kQUNzVB3szRcShrV0
L5UdItdZ6mCDTyo2AraTytZRNM7CfkX2Lw7aW00GemRZPhRG9F87bIJGnA5+NmJUs0MgIwJAl7+b
TuYotMVT9ku4fyzd4/GKklV09EAhGIkv+9UdEpJI0lfgTBFlcdateqdF4ZMQ3Kz7EstgssBXM8k8
zzC0SoSqZgfM3ovp6/XmvSSUJQd7Hrb4N0Q+H2cGJflnsWXzJh7PVFQWWs/EDodYku8UGbDXHtSg
A6KzrGE7R4f4Vd69OMPFZnspeqXHC28cawyXoceFR7FF9uKsfJeEqLB7AE+cngu18Zi0eUWJajqw
32v2Ncoe5e5gay1vCZnUYA482DL+YWDWOD9PZQmQ2v6l72fdlf4VvUghguAsVHAgpUBllVWZL244
aBNZLhSjOF/ALivjrMDPXnzNTZTjcYf4h+9dQQsI9bgb+KMAz0bIujzguHQSHDxEYKVhFEr386D4
2bxHUh8LUvHthlSr2lj0Az6GqszbuunoPZ1WAEtXYYpMdriUlPbx8bOSGT8pHnZb8da+j+bm4dUl
ZG+hUSwbcvR1N68nzsBE6bONMaZKmFxtOioDVk0CmF74qHkemZzrSqQBp6g80e/1PEvGukXrv3Xj
rYrPiEW3J9fOSYD9c+81ETeOtlDk7tL687Ny5LIxlGJal3Ry5O23Q0D6yMPJDF1vdvOiHAAoC8kR
p1/UTc3W4ikG9jF4wCsCw1jU46HINfzbh43cZpfmzyB6tEuI1Aqu93LUQBfHKnXw0C7atvFkF5uJ
R7k8ksPxzwPQRhrM+IuvKYr+4WuShMIluzhPxt+F9Er0X8J7Z72Uw3xZTAgCdTUv2D4WuFFXlwO6
mLbdlFEPecALNa84XFd0gJbYx9qo5ruMWSivb70H3QbwZ4tJlIBqk1eBXQsF/sEnYMK+omFko8p7
LTUhAeH+uKj6z0gRCGl1+Ns2TDzsRkLMfJi820PQ45+/QBk5trIkrnIR0KN3bZZYS1r2OH2akW6z
UZqbKgUxvzgVtUrzzLebNyIYP/iIQqMM+Kgm/Bij0urRMq+k6LmdnxZDFeuXpD8XA5AkFMUjuMsh
WzbdL1JgyECFQiromlt/C+Vp8j09zkivkRpK+HCJ1az3G3n6Bjs9dt/BEiw00QeESfFAzJMoXnow
DQnTxL4SvYnFVK0BQ1bptO8fNPPMvQVZqKsWtDlkVacaswAZLkoFXtnq3Uvea5vPgQIS0jd6OC/u
cHatQC4JkevZRga3HllCdD4ugyzAnCsyLnb5KDUJKyVsPmHdCxeR0+l+Ptglpifk47aJvtD35/SB
4A3KQIninQC/j6S0lCXrWn9cWDwDCrjrX/NoIEo+DvezQARH8BdPApxPm+Clq4iYV+OBcxIiA4ty
JDgKq1+/bBo54Ppskjb9gFKr+Due4QoVBTJ7VFtUYiZ3QmKABl27zlBm5jkgT0nJtheXl/HzPTO3
aY6kCQLMCxX2qCbq0cjIkMlGKDP01g7SzrD4rQJzj30CZB8eIvjHQn0kjw0AgD0/ZTte2hL37jta
zCfVFEiUZyqnuhEaCgq+VhX4XTEKPavQf6mfNzj1eH2UA2m2SccsI1G2c81gMEwKM+FmhaxkN9f9
ilZLX3VLCC806iGIQhea9QUB/tCE3Po66jAm5i0iQrEN3JyAxA11sEhtd044JGlw5wK32Sp7QhXj
2Z8jKlbBwv1SBGQGqgNuMLU2DAm/rS+KdVF1oijALYgUT5M50H8HXX4J9gMOWv2bJ7botfggHxHW
b/w+tTqSdQEn6lsLez/WzfFTSSYKXZSreiQjb141svkUHtCS2rwzkeTMeA2sd7hh4+PtNiuZWHs9
Fx1iCzmWN6Tx8ruvlTiHeq5bPSa5dEWLMBB4/fJj+7Z9kkJbHNX96CvNXXVFeYy90REsU59Be6KF
KX8Bw7lFFEaZTaOYA1HweE5CDi0U/ccZ7EORBhVmvYYWlJxSx+w5IQifizuSm9AkZNaSwC6SsK4U
Wk8ZIjznrvejao8bsniUVRejJWOc6WafjtKVZIQjeIrLtoKD7ZNBdGYlWc4txqz481OmDi2mmWIg
b9umNFKbPsN81fqOrV6+HgZcnnVmUMJi50r8CQhzZBxuTpQUqkWR0HbkGz6zD+PPaxNtUyyNH7y0
z0C+x7SQ7mNVEgeh0wsm8H2V8anrS0ZMg3Kb5YvleVM+IOD/4fdYzA/jEs+EW8AeNHIz6ePfAFI8
zoOXt+p2lw8DQQ3zQZSrR1y6nVleGxh5em/0fxLlTrrHt7dQD/D0/AD8QHFRL9w2/r/Z81MSReVL
c1NmCS4qy3Bw5l35Knh08e+I31Pqw7VOc7IrrUYfJw7UUS68NIAn6t0p4h/0XPalJ3kqezwesklI
+4ROSWOFyPr166iyqbygH+mHaUMDQ9Dg/ewkn9fE+NxzXctBgGE4jnsRPGguPQoi6TU/rJpwTEnE
XM/yhka1WgQAZd5bETLxpY8KdH8fAK4FnxMTj8vNS1n6EqdpdcJngDlkMSOJzqCyUmyErPBeN0Zw
nd+7M5gC7UeKzsND6HrGqp9rWpRIisrfZCf7jpOn4lrOj4dn+ko6m1F8d3RmFv1C2xiOWKnl+qBM
4uRiWsjU6PCe2qjQQzHoUUaLv6vCwqlHSICNRasTwtBD4uwF5fNI4WqD3z9IONjCtB2uEc2z/Hgw
MPKO3a/M2w/mpMhxYjMkZ435LjUGh1aDN6re0/WvdJtUBHV86QT4RpkBixH/9NOo5Ne1tSg2f82g
+wCgyYnM6p5KU/ZoYw54Uxm3K2yhRBFL561UCh2GlSOnt92ueZp17oKJiyswa0KWl8Efkm5M6InY
Z9YlpS4FHDibP7k8fhH2gnQVG8EZGFdeu2B73WxfaV+MqaXe+5kf3gr5wkcPy8kWIBw/SnPnYYPE
DHo+iSeB/pj41C7XoG0t+egtTqzoFkdQS0Q7uvRiOYwAqzQA9BNl8l5lrdurs/gN05ec61LVfTkf
B72NHRQEtsEac9lodpJBPpvK20/jPb2UuhYOaZnF9ZuF/198/LF1xwA8IO6D3wImSFGTtQHDtige
HGd1VvkjH7v2i7dwbFBRFw9TRFSwVD02oljwC2nyaEBzNSAC92IBAF3RLA+TzzohH6A4NTcBOppQ
U7Cp6v3baV7EhtrNow6PKGnmTXc8DpwrntzT3/S/okmsll4v9CL4Q3gHZ7WHyis01o+XeG8KOMUO
YDoGhSt/bwpzsN7h8jweFzKkmi6dUeVMCBgnKqAe6FqRnA4xYv3WSmVcyONu2/i3rFxZtgUy1SXX
4Ny9ScL5br8n8I2W0xr5EsMmkt5RJOLeLs/2gUC7/qSv49oft0ZHlXdecJOxilh88rjABSS1G9x7
WnITL/oq/b64jwU5L2yx9kQEfe81HoQ2l7W0gggH2R0/6GDO5lsJX6ZHP3G5JQGU9RQovj/6PeP7
jYZoYqtf3Sn76896YJMUs7OZad9teqm1Mq0EP1/uQQ8vCeX18pqezhzGEMc6APcfdln/nmHgwCy9
fGzsyA+enGtQsqpejjoLgZBe6ZqbU5km00tOglnN9R45YLMwDBbAsf/chiNKKKXtbp+9OIwxZJhk
5xpJg+X5LiiHnnW69MGXScontlDNjyEtI5NQ0SCHTtYhAeTJu8z6/KbTdvdKOnuf853zOS2XCVeQ
Wc5ptmx2LWmC8RIDEe15cKOJRkXqvpHBqBgHvG1ItVSmg5GaTR2dcyOuzhM7VFPP4DqUoG5S1ytK
xulY0DFX8wAC+tlSN6lajrDgheIfZywCrNzBTOsMROHZFSsY8Y2xZ6KIReD4divh9AlXkubT0x96
RE0oiFlywe0lhvN6W4ApRFNmup0JAlEaTKxVSTu7kNeFZ+Y0ro3B5Y+Y7W/FySQGky8ilr3lAcrq
pSmEEfIDPPuar2lMnOAWgsuX74tAg4PimbJqI5E/vjbTfxZae/JDVMYfCo4C0ltEEXJPNBbJ+8Te
EA1OOTtFthOnHL0WW8OuHBb5Hv/+0Rx+VIAlUxhvaVKFkxtfrq9CdzQCSoOnsyOwF1DUSxjT6Ytt
8UokE4S3wsnMjjvarSwhKRdH9Tdbcs6LlR07T6lPcfGrgs+RWe85oYPKEa9vtxtQzg8EMIRYqKe3
jcqF8eRQAR2mEplfeoSnkhGvTyTsXsL+TajOfXBkIELglzC+rKYfZBg+KUU/qWD1DFG+GL2JJW7a
aii0JeMJox54ynafTZ+vMzgdxhYBcN6WbFNZ9AJwvdBTTw7d1yiXcRiHXgH6B+gu+W+Fa5s2Shf8
gHW3Xp5RrVfoNiEM9itQ/ttLqBPjKBhAftAhjCjVE5qD61o/MbZGg1JCUtKPUQi3qJm103WyQw9d
Yh5z1WUT4RI49IsUzK46rCkKB9Y1e5zZYtedMCRCjkW5i/U5KcNX5ctdFRgC9TEt9VOvLzpTwAdv
M+at9feoz6OhX7Kb0OwLzgAy9yNBNLKxyUzbQXv6CT18yVOeSftS6nFgIKtl/a0YipgBe/miLbkL
fsrDsrXmIjofAVhxWOtOwPK8+DD64MIKKwNtuvf+mA6j/4E6BLIgaXPPTcFZT3S2hVCHfkkPj8CL
oavjTR97DmXAOwOnquLmAWxdNi1WpjiPakkgFksktyBbOleOckCMBGac+xOIocArDxlNon7rTUO7
Q5JSUOVssUJSNmBTwXLQr0DJRhABLV7utmr+XLipWlWQxUxoJCOD2q1/rNNaoO/W4f00gYsKe2FN
xii3bI9KqpybEoRRAH69Q2D0JPp42hwz41s7p+23hNAOtDroakAWIZk5br+rx7KCyxua1iOsmmgV
mZm/Bnf7/rJEmOQoIJaYrOL2oFrZwRs0b0dqN4zMvyfLz7EXn+JFBNYDSaSzMykcxR6esr4t7eHN
+YAIur0VFJVvZ8wH91gM5sWDS30xOm1h9ggGooB9iNtl7JfmyGdl9osfAGPY+JnZeL0Cjqd/hmKI
P8M46rgapWrqjlFmHibAjGKHqezs/djQzqOCSCt2BZsQ8yOZyT0eZFgomLQ66r3jBYBzRMPWdJrR
jvrLP5P3Hm+rEzctJBZCiwQcCH9C2gaUVOZ5VPHIXcpvYCBH5IzP5tFX/DcnJBH8cYe8bGv4ZNY+
dzlb8eUEr95fpBRWJ5XF0q+H8IH7Ob2RvD1bAyG9q6ZhojN5WqScSoFPWZ9IAtbNUsaknq3J4KuY
ky+R+hfNnuV5j01sNMpFJUQjMsB0KQCJtJYC17xMUJgkVHVX9M1VJWrEvrvVd1d0gHf1HZ3jR3D2
s3pFbElG2vc8yGK4pKftHF6JyBuXMbUpRkZN1vh/R6bJXUR6fk5knUi5ugCLDvKa+RknprpMB6jX
G0eI+C1GWyOgJojGxKGFQSBRedLV4JaKBDh6w4jj+mdvZA8TReCrwBG8Keq+C1pGkfgJYnt2maYZ
aMtukGiNlywg0S19n1oC87f4kIk6SP8A7E8xE665YygnHDFlKHrb24If3yqSvzgdWefm5kKDy+nE
5qzf+nBlG2hc6QGitDIyDQo1YkIOENRXmUMAM50kS/k9i8aEU13RCugsPUbiWKBEiXDm+zDmtx77
HlSH8bBWzk8gvo8ThSps5LWg1HILkjxjLkTrshEw3KSFPoqButkjeJ/bPFtefGfgrylCBmBTS89d
w3kSPCs2lXZRPeexbQMqyt4R8KBfzIgQY55PEjq+ubdBz/wVNbxD8PnNBkiSPnndRHyLlYxfKeYt
iLwY83z3772sAcwCXMt2i2d8MvFyvd802QMhtPKQD8OMJG0Bjp939tL0oSN/qGwney+SZEJlaMQJ
d0/bCnP0cccnPoBvP4DNZDduIBpP8rNmNaohdsBPcmKPLCRuscG4nj91mt8IG7le+cNgyAf0MRb3
eJa39yTVslLSe0UwPd6C3IVVLz/8x5y3+shrVKxxO1XBLewwBbXhskP6xc8fEBjv2F8PWpBj3qzE
0NJb1mv8AtyrI/VyMFpDyTNpuMHnl28pWTviXTDXN2lvU62YHySUdZf4jDVYxE2bCvdNeuVF0dvU
R7K8D0+rxJ+bUeHDGQoqqJm9g1N4wJmwrJpTqFHLxIXdOOnRYTYB5L27uOmW/CsB4fSlE0e+Z/gY
5fyzjzuB4aPXKZ1oICt9Il2RUqGtH4vwQs04QIhFKvjCA+q3RXux4O828Nwzwxa8VkGwFsuZpmsy
kVzISqGyNBQyyt0t2J31aSmBQsznEwzBpdpd5ilMhHbbYHbpBXbxARJSTG5KKtI8moY9vfDvA0f0
wrp5aSBXQefLQF9MiPj2U4gTUYtZqV09QOYIIiFm2/DDJX/H4yScjFvkrvCiRLJiAGO5f3a88Re3
KbRa8pZsJa+83H4k+zSsGHlrBvpAq3sM2SHkxMTcqUknuHCl7aiTcb7dTYSQNp/fbAp0ysdD3UPM
pOGwmFos6GEJn/Qf5NVcZKktmELPFDeHEEcmCgv4/EhuRw80WtFnBD1FO+hu2Q7BxhdWqUPDO/B8
tpHv8tBVOKs+cPyMpMmoJIeQ4E3G20Df2uaihg1ct8ojid32eZSqCqZhKDOBzTNJKWhjlXcr0JOQ
JKcECvRTqusr8isB/0W2yQf6grEgIb0wNCt5vIZ00bM+J3TJtgPZvJbi4GKtM3zEz62xmzT/ci0+
pE4LzTvFWomuWIFhyS3C8nTeW1LEpdSATBtKjarAexiToSvUGU2qwb+JZqpVYk2VLZtY6+R5m/lH
GVNlw8rt+w6G5RFAAYzdxjvdIcK2oMwmDIm1iMXZSkQtCbr92wFAtwRf1OwTYiGp+ZiVHXHr+x2h
vlcZmgyX1nGM2FgJnAL7UqOYmL3MvNxtaa6oTAxxmEIfcn2PaWcAouWkxLjq/VkB1Ul4B9IuWjB6
2vGbKG1L2O7DSMZ1VUnGj7SdXwXv4+CEmd872KFbRyrw6LMWnBvui4KnevAC1iYrw5Q8D32F/axw
twSeurX9MRJ9XorsqJug2Nn911QPw+Z3XdlZG8x/ZgPKz8VuY+XBlRoAQxfMgWGRlzOKfchuTZ/H
of2o1uKevQoIIA9PacBxMPmgeILpvCgigwXoOicmoYk71FLnS4rR8HJh6vMJhuvu6KS9fGWWat+W
PVOVPVPQPAps/yCI7N8CQAopmifIT/AgoV1CWnh9eeNWibY3n7LwqcjJxRwLQS9lJpwNI++CSHsL
Z8krXJkEaHnwFhnEi/iSdryCBrwp8mmOK4CiCuUSqyP0EdCwt3RWxHAsYb/KsT6zX1NKSyBEAgfT
sKjvijkYwsL9e38uoafjkuqG/UmP1YOOvJBFwhae3X9cOSoJ9mVbLnSDRHlh3TsOJ8WJjkWGXcd7
lnGIiemKp6ZJkiK3UZuCKxtoVjiEIs9nv7wyZduoYTVhldY0R0jhegJp7/kKiilRbswhen4+mOWk
R69czE+96FfKBbcBCmu94pb8QhNkcQoGKu60l8dbw+HuhoxldY5IijsZJ6sTO3Rr+Dco5dK35khW
Paq+kchrzdSopMKiyvEruOCRVvDPxXGv98OxBxZmgLhj76CHnQtCFyoI6WYatiCVmCRH1klxizt7
N+gAyxR71EGsnV+MUebRUTQn+pnvHYTWT2pPWv2//Nwf5t4+oOR1jlL4XqNsKjCJ9oooTamMtMoR
28VvFUeohnAdhkCxmllqRysVVdobaCuF7EX91Lh+Zr+P8Ip+7XDPN+B0oIH1OuK+SYG7o4wHIawS
0gFoVwsxG8uv3jYvG2oZjsnNki3CRfYxvl/NnzZE9TzrlPc5ElKoLes1Oi3zO/sNRoamK4VhRqJT
oMPx07KH8odpAkTrbb46/M0w16Ft3CkI4VT4O13LcA4JTyn+xz3BGbw5/74dpsTk4Hp65/2Wh1K5
ogerFFMetaFKnX4Pkq8xLDV9ZVWvjH95TSermA5yTv++cLK3AcB0gBfakKx8tVluutJAXFhO1VEZ
AzimccVkiIp/yEYZc3aXFVI4H/mqV8FGlbLL7fhtns81VL+MqYRNGjIZaHkJFuNOgcm/bRRX1D4g
CB3vtZFN/A79n+OgMvK7JwSV8vZdH/viHwLw8r0V/NVQvHf+V7gs7QvxGMuPckIQlErsteMpO3G5
GsQnCoJ/YWZ1jkysmVxuIIQw96eat/dqWbGWBS+nrjaEf8paGxDC3XSahRbXJpaZ3sxZFCdScAMV
gQWkZz0SNMOiRBZ6NcHzQ1lvrYdnz8FYayfGfBuI8IZ6xk5ux5ugZ/2HKlLmPFAbglHGdGshivKF
R7VeglfCX8B4ymsCcQokgEU8N3QoqXxWRa699BUyff8WpC8y/4xmjkirFO9rnf9mPd/rgIc/oJAR
qFIVbU80BtWYzo2Dn9gSNUwJzg5+Fl795MF28UNEGJx97zBQK2+oaKp9GyvcY5QItJfGKFtNvw7N
hii2Dem+BL1c/EUWPN/G0uKpH0EkwJ/g/BEqrMSiJW2gZfYvDkrhj6KykvnUmGca8Xw/AxhKSqOb
HnWMjlY5lCZAyYN0skmZlm6OSi82AQE4p3AoJC+YfM3X/DbBvPdg7LjdhWpfCUgWxfYS739Ba7Zy
reptZxjPDJ9hyerWDY8FmSKSXXeQuO8milOmCGJavfapNP6EZVmtndUdKn6K5+ZOVmtXIWlq6qFv
27kRBx456qIHDRgQqqZ+t7NtuMWqxEoaRbue/1RjLgGBCehuTJoFK0zA0a2tWY7JqXfaH2qLqdL4
8HGR3eQID19X4vxSDOfWLT+2tHWAn4NPEiEW601A8PlDAPc8zUWaQmSWOo8LiPb7HjJHjAe3+HPt
8unnbYFdLANliBHx5PYi9HS2lDo8kuIJMAw0xAhsdj2/9vAUABpEiZYrJSlUl3LL62OZxkCI0394
n+atR+qxKsjkYI3WVLrIuqQUIqyBqoIQvVcKQJwfywy/gGF8Otdk/K56GWQSen+4QjE9XkFA2HxT
3oDNDl0Eg2FmHvMc03Tst9WQ4ty4PWJblKTqCGYBIjQ+bqqSZK7vV1w6Pxdyw8N6feYN11zQV+A9
5Voujz489lKDsC9yVCsJDxzjsVcQLFmb+xPnh/SqZbLVMhDu9sthHey3ryLgepKkOfZIb+D2GL40
I568ZiCjxZM0srqNjdISt0Y4+e2D8pERajVm06obCYELfWx4cAc2AFSGUapNlKWGE+M9G5OR5NfJ
pz0RFv5UCvfffLhRvfzIH3MYcKbzcDqI+l9hrPpDYnZVJ+Xm336BVrDzCDcBYqttbQXdi3jiDev4
u2LxsgDp4E1amweJow/y286reQlxg5IaCWcKyRAq6C+BwconrhpRCFBM8T0gllwrQ/NUNGjRlyy0
tfDoYHJWKivtI0t0FEpRIiVtSk66xp8zk9gBqMmN4SxrWoot/bIpm5msH4aloOSKrl45c4WDLcF7
3bd1LY1raGmAMG2wwTVzAyroYsigls228dw7zkIVkhuHTSYgm8AvnFTgjj94zc5D5ngf6nH8OHNi
FonlltQe+CWgPaK9k99am8XUId5SE8B4h9X7h2TTLHw/GvESMJJ9QiixhmXq1nzWh9B4tVqhhq5Y
RdWGPDevvo/vyek3TvL7fqxygwWt8jHVBLBjvszBuIBmGH/ASEwRYn5MiLtMsx6ObkHKCQpzwJAl
3b/IpSGZ/g45tHyEj0V6EGi2mdyQ1+J9BiXrn149FHuLiR1IDjYKT7FSe91mJdMVqiWZjjyzZsFA
IOUMsx9k8auXtoCP04VbCLROR6Fc5yDkBymZiGAiIWdcEINMnT83pZBpsz1MVTvudjhreM1Og3aS
WP/8rPd0unBPMBaupFgdqM5fuLi2UgD707j8BAkXXUHisk0NUIr3zaTm+hdmwlRan/FuzuvKk+QP
ClI3kRQbrqlkUQDVF7hQ0SFcd+9BEpDJgE6ywOoDpO20eTmRyRdHNXz/j1ImR2gsGrMtAuJP1kjx
VERNfk9Z5NCrjrsAqMPvEPCvtvlN3IaPMYLY2j3jTZMuddcwHJREKFpnwu2GhxS9/PtKW6Vbvdzc
lTAvjOdnEmeLfBqxEhNtpz79G3ftNfP0ARLYtFLp7XG85GXWrUOj+k62gIeA3wRpZ23EEH0HEnL1
wPFG0rZYK7y4YEQlRGtjsrLohAY5oli/zVgkbieV6nCAZ06SmjiKaclNsMVyFkAvYtDsmVm8oo6n
LD6EozyU6VX7NgxQt/rLiDdjWRlV3SjJ4Ik1sw/z0hpbZ0dmVrMqJrqq89j2Vtt9vLjgQzvcE0re
BsimRDXC3eMNDshpV7bRLMHLMm6O+K6BQB9Aa+V9orw4t83Xrz/rzPbTjTLeELktJcBf5ZVARo3x
/B8SWj2xU7g22SzwkjGgn2GXWHX3pFoxeDmWbsE7+byCYZlErJusxVNOsGTSSA3+at/BjeTt10Lh
shHjwcmAJz7fDMfmPB+FsNPFKm1eKe2+sx/xx7mgS7l2zv2+XoAxQgblbm811z10MIKm9RP5Kf7k
SvLoGrM5uEpANknG6vnOQ8R9BF6U2dUWA3khONUJ9WyT+AsEXewZ7MvvutMvAsOrWG5Wng7TcmoH
EwQwg03NaZAa6jxy951vPO0/pPkWDINie9idbqPhCma3k1qHqfSmtQGQlwYwaTBH65YtxnoFPo2Y
jJgOv2ClP1bW6uzI/vuyAFL/zaMIEMC13thwRsg0Rxa4NaKtaVHP2LgWxhzKhvAuZu52yEq3ndG3
5/BoR34kgY/yOTXfERLp2SodaGtatf2IDCyjgclU2gSTHAhZDZNnWV+PIKisVvLEcWrEBgSt7Un+
Zxop7J1EvpA0/+PjuvOPUe27hBC11pFOfxBuCbl/JSg53FnVP1RbxbuC9zkGY1/IbKzx5qFraLih
iPCw8BtGqOndNH+Ff+uVETWt0n52C84mJ4+25B39m4+y0Zxmd52shQCb/0nl7JkEjTLrOtGsePJu
OmJx/kn3yBsMOChsGY9IrM+VWw7xR40dqz0Dx1uRQU1Qa872KPBXsRON68Txu8haAqm9t0raAjhp
IXe/Da9r+2+JU5/xGS/Huv2XkKtErXh9t1ekGzNmESk/ASorOMz60oqJr/fG5AhrSG7cWlMdGNqu
cndNbftIgsOrJxoiSmWYMqn8FwWHJWFcW1JTz8iPJe3Lue2MLIAXM3k9y/jCgwaTIv/2pbDVfD9U
8zYif3mLZbwFl88X4uc1ck15AYvRByekwsSexjJqWwYC6/GDUZ3ouiYe548VrRtOxdo6wRjz1Gya
FE/AE8dDjUe9lBm0HJiRLyLujs+oUYVBXXg9/C0pS05NCZcTQCMpaxjunEtWmHmnGxm4iB5IMbit
7tFUrI9i8xcJqz/kAWIfNbKoK1TxhLcszzqoPq7t5LJMrBtzdLHBOhHvtrZufa8PX4OyjNbxIUx/
p1Cb71Yu3dU7U9p06tiZ4S18hXTC2gq2t5xOivF8kNoZb2SHdzZBoFah2BMoKJIBu8z/pXne2WoE
5HlO7XsONQ6NiD9lc4XAL7MoxGJfisVdgMpzTvyJfRq+01YOn5hUuQJ/dLxj72mBWNEtxnSQAnM/
mn9lsm/omi2w4cPtktsrglhtkkmvf9GOCVhmyd+9FFmr9RHWl8+436ajqoi1+gldARnlCSQAxRcn
9QBa66fBDbRh13YmbQnkcnZVF54uej82UC8mWZ9jVsXWGdfncZGjTZ5BW3cIfNPAaX3ibH5ytZeQ
dtcqZ/Pw9NaBEuucYBPdyzSD72tzUS5SaNx3LRyk8YkOI58HsOCPcckZmxIWYfrHc5JI8FUgnmTN
mWXAzxJEPTvAd9T7vE/NM/yO5G8WA7OfLQeRCXD7r8bPBq+8wiUOgKEoyIbaQ0/oO4vEl/8hgPqS
yeeWzgoIVgru0hA8Go0qD6QVgDTVLvDb07EvUTbmtmUAt5scWyR+lN9FX1UyqgxBNdMlIMn60pIo
R0jA2ZVJYLne+J3+2tRTa4EIFVKbiqJq+9MgSRLsRD+eD/2XXHdytjnHc6RbPVrDeNc+Tig3OqxW
aEOaWnSpl9d1UWe//8KYvloF+4cjhGwrArbvBhiKlTohaTyWm+h85BiV58XNf9rodaWwmbuK1fdq
jhRF3psNOTP+UnnpW8QkQlzQnhMpRsDWuGA86aovl+J40oWcyTS/EQiUi1DDFXKcV7ntTnT7Nxf9
Ysr7q6zDkvpUx7E+u+ececifywH7mULk6Q38uIppEEJBPkun3VD/svSKyl5NqYJlMZwQOPp4eMuP
c4n8NJUTPDCgZGchEVT7V/000IH5TMLBn0zssD3m/g3UytviHh3ceZ0zgKQGJAMqCMAkspuDuGYo
AptvOf6jIevxtq33n1hd7pxFcpqLX8BEIZsVg/xSzNIc4dBF0Y6ewxtCQlV+MbNHGYJVIOvqZq1m
1XJ+UbAx+6AD0pqSYrwwYmDkIsndhzHVT34dsAQsMxsgfFolZas13mXwF+bSXEqns6NMVImLsxev
1rtjEMv4XG+RehjM8rELuSu6mP1pYQxJU5PG6vnOA4CTbvJtiGi6HXJO7Jfdek0hRzq76Lycdj2H
wjaAPt2yLHv92UfoWLPTNfeAouDNXQvBlaK641R+ZFFmLiJIxhvCr3upIOgn/XzY0CUqpQllKQg/
irGbFloaZv5ymBXcsPVJiNdLkIIO7oNMdSt6l+vEkPDPkJPfqW7CcR3h3whb3kQzDRvoLRFA5DY6
joCjJmxIzEr4mJG3HqlSlxOnzdv/tzTzsMKvs3CYbXIG9qkrXaxVZ67Lfeh6GWYBYfTMvi1YH0Dd
CFgie5BZ1aNMgrDauc5//LHxnjHWS2msJI1QhFjMEHXnJjB1ATEsOozO0Ovo5OK0rEdAmZHSr7cy
Tc83oTr2mCbg55Dc+e3KzT1zeTaSHc0QHwHJ4YcXr8YOndOOJ2WWUR2hoIptt/6yzhhtASrHIgwh
UeKt8E7kssHzi8AmbpAVGy48zTJtMIardqKuS6Con/819aHrX43JxCVEgPMXxxQjEbmA35gUv/ez
gWs77/ODETsWCICEuDUJlM2TnO38IE+csf5jSC0fBysk4RF/A/4hUZ3mZ023+7OSQQzsaAa620UJ
g4HuNOfRnXWrKjyRN9jePTjr3A4eJnCGYDhrKUVIhVsq97578OsYI3TU1we2mmZ4Ycmz+GG/WSVa
y1pvLGTr9wsn+uoB+f+rnjIDE5v65CInk2+gkMCWkk7Wa6gOTFMaT620doJhv2VGWSa3HJLpnLhg
zKBzr49/YHSGdMy0xwBRXmeeiTyfpSw5beMqnoQORCy92HBm7gQXClZIOdRC+aePqeUPpCVHO+CS
ZUEwFvmscU1/LiNftprZP9gxfRCLwP5GR3J5NH/Hp/fR7RGGOLTtsQdWnNpZjWWDtpYFDhoZ5oia
HnEP2ydkn7cZNvdzBjGku8Pm5kNLtVk1R5DG47EMBTG6wukwwe9FLuTqeKsGLuCIgUalnMzZLzPP
NFZzevh8aGo3bsBucGJfCBmPdEq3jEdhpUZfbVuwI8zbn0f+P44BqD0qyYohhduWbSqmGsrgT8lH
hDSTM/2MftvgEwBmNhNtmDd75QcSeZRQNWECOa3PI7Df2Lr18D4RLfMTTfhZ2g0VLsZz0h1Cahbn
zWK1zcV+sfUjEL+PRf2A2kcHktQ/Icm1win9EJPvP+HkSd8N1+yWKPKwPE+It2EEHE0PrZL7gEzn
reJNdV63NaN1CkMv8OTEWUuC0NaW6STtE9jwfhmKA1ed883/a5fNLj7Yc5c7+UMSkQ417s52yScH
a2IumOqRvQoAXkdgrXvgI0Qwg36I4MEGG9kP6kJ4yms/d9b44uFSlTK6nMDv5I1n8gZP7VTE4+wX
VqJEC8z9CQA8b0F1VqDJ6YRiPoo+LIJjIUPF1q0p+ktDqUHMJu1FUkdnDploQy8u8pUn0Y6kJmAc
5RhQeAGwpYUMkVtxVJ49Ws5zSZgaNMqdjYGhAMy8jRbkHcIXBpNToklc9N8+QAKSk7ANCxd+Yp77
w+BVwAQSaZSZkSgtwWyOd+fe7ttpAOkwaIB4WWLhJ/9ZvCVM/++KWE7pb6SxV4KVx30gPwzsBkAy
iXMYg/d8QUbaToaWK8bau1YVYUTwfiY4CyPkSmHB6ViqOOYLEU5+/qxUzCjxmIAwCxPC2APvHsLm
oNQ+gdA5ly6FD3YOLAVCafw6V+nDJnCryh4T0T/HCOyf39gKpE2U+WgeR/oUF1B/7tCGkKPDsKd/
DOu6J3gMt9/LR0dx8PKG/jXWK5wsVJNQ9KdLGO56Le6wgjWCNU5NDugllY3N7kvIBBreYOlmbE/L
b/f71k2XCKm/OjlJgCcS2gX4FpL4+vI8JsKSRxbg/ORc+piIwJ0AxwuoMFEeH1laxvG4b3Vuf/OY
jdcvpYbFTICzns/bWYfNMjgBvkIqv9nz0uPs02Ku/jNV3IFaqYaARiEte4ZQUfjU3+jWqesl+JG0
pdtDmA5qj7/r+XV2olJMTh2Rdm/DY8sohP6MYoIsdPYPZSLmHqehUlcihg95HI7H9HLwTSvTsR6z
/b54JLPx6qkrzvmqPTOZTBVDFp/gDRh+zekSIDenMt+QaH9Sboozxi9v7YMasM8W/sQJT2MlOpeS
0sU2hxEwYdtvthDVAb4TFmqNtTxcDRqfJb8KoYgTrBmKGj8bF9HHmkCeRQ1iBycZ2YS6f0JQhycl
pdNI3yZ5+ws3YHdUxDU1eY+2mjOUINRoh8XL0NmVm2cMNpcQbXORiHsQPJqxyMgaySTE2U2MkwSy
huMSkkScg3kxT6dVtf+JitbItB8Ev2y3Z2ZDlaexGOqremUmW11vpdvaUplSex/sale/E/0YCIyR
wfSQqYVMN8E+nEGxxGH8VvUBgaG4vAVWfbBEdRuXInjdX73EvBwp+louykMu2nkItGctmR0ZBh90
MrFzpUWzved4NJpjTfLPVtNH1xW77NGTN8e0l8BzvL9Lee3NgqQuf+1gLTE3FbZM8ECoFQy79NBC
wrGf3aVR3H/bn2VozvzK0Q0KFP4OL+Tf1lVH7nnYDqzxV2R4QrsMgSq2j4coyLyqibQEqZZdJjKl
vUkEaXJAsrW6Ie3cKHp3MBsrqj4vPVGXnhleBsTMLf6CP/GBRDfyicqgjpUY2/7ttTxYCbDfLnmK
WM/ydpI6tzBSytEiqrr6wATd0GUnLiITw18d1ymWavxWFq3G2zmCBgWzlotPTlmAalYb7syGRaY2
ZtjVFL/IJvdeFfC87R0Z9LTeuzDMcXlvvNTRwTE2KCAc8xkH+Tc1/SpwkuH6roOoDMoCAhI7/znz
AAHRvFWROGzadK468IYyBqDIMpKF6FvYwI1JplPHQjoNwGJB4ZGR71zVbllddFcmCyySxAynBo+G
iSn9LVxOvXHnqlMJvx0tZ9arXnZS2gPqI4vFkh7gYJXszQYNnqTF2Fe9wXdoeJt7pURrKdTOsAVJ
JTOXqMcdckAMp1mh7IizxiyZAI/jpCuQwFvvldVk3pNFqhF5/UE8LPZoBb8NTfmEHkXewf5pBpM2
Lugh3qo36j/fNCjtVy4mAGT26Y9seeOcNHP9ZrBdtZda22/kVqg2ZV32dZs8OlHryOVf51atH5ZD
QdvRu986VD5BNvVeWhTFiocVGJNgfyhNQYxH6Q0WD5K1lHEr7LcADG7BFsCmKn2P4P9VzjTgL/Kj
QhvQ4/AVAmxJEkXT/8qWXuw1LbnxtdqGPQbERDP8f3jEGz6XpQhyvHRqWELdSWFLWooG8h9VHTf8
2jILBxBVMicJTA72FrhkUNTEYNvwbbFQjK+au40NO1Xh0HmgaSX5QDhVArtXEz95QCySdK01oRJh
vRChcrLO/J7VbLUdQiubTcAnbv4HfG97Qp/3jSpys/Copma6Y5TdUns+jsmgxY44KW2GvUyqThEK
Q8CpQf3CFdtvXc6X0E430f8PFz2bFXYEtPD6gpsXb5v0KpDT/tSXVjBDIZij3aZN5+q1268yywxw
VQ3pCaZ4QzbP6csIA7V2xEc1ur3LE1i6rtJ3nXyT93VKmkmzWovGY2lTnspLhO0peiGjYgyD/uLN
+AvaQFror851AtOi4AgxPkw0eAoRDA8L0ngA2t/CAONz3mC+cJcn5AnvCKfO8P4uahPXR2nf7u9M
XiQUvcnWZB0/Saor6p5dJp5fS65hY4/n/y0o+YTH5ODa7QRXL907CkHIRYFLAJZvjb7c6eflyooq
AJLyrhBGcxrzXqoWJTb3nN9CcJz5F6xHr2RfbiDGA6qx4+tYDdejbRkDVmSBSD6B+RrwwfgkYTlE
OmmlJZ3Y2HGt5fj5YIAmYIQSOsn79qc0fi95FSDn2GLmnbf8UnSmO+uMGh6s9UZ9CT7JfRstS7P+
kZcuMyAE5bDIvDhN7ZaCcnQv8ox/79sR95V67ximfQoUECbYodvCZ9pOTQXV+uNaRzuf2ZThunCH
OSqm2zRCe8xONsVqCH/RK56LF+VEz+bCUi+78s4pMZZ8vsGNGH8LyQwBspSdgrfhbRCiAk1wEuAg
lBbqMQeQzeNfUjzRUfdUBVgjVtIXy+z0bEhFKNwhlCeoXG0Q2+qm6mA25EkfDzl+CfNgE46OPTlb
bFrKcEmLlifUAlII+MoRB87GgjTsYJzFFjauPOvFwOviEG/sDwYy2R5V8hJrND7txTvMXfM5/Pgg
nzpSDQdLs7XOEbhdJjJHYPt9wT4o+RuEMR3hafTzr9EEuBDbtIhpTYEqEG1eS9rMunEfGIsbNJ7D
u1IDOIGP4kyfyIUmG5SscFoibwYuBNoaUZ0gBe8GZqlHNYYrxcHF17suqUiXlu7SdDxPRu1HXnN1
/NnyPND1mi7v+VS7BuoYYv0wS9WQ0Nt0cJfQtU8ggzmOuETpgXvwlJXPGz7ESHJQwVaUC5rxCqt7
jpe+yyUxXQuJG46s57VyLjsIOZWPhA2eEloBt7/DKufwgJ4PfFUHMZWk1GRhU/MB8CxaOxlIIhuo
UHJEXLjWXJGt4vT2D+lBAfWZglN+u13hd8SLVjKwuqZRoqsRHoq76dQ6sf+vl2EBlTVAk0s4p9hV
ZI3o8MsoQXuO9w7hJC5cjTirdRfpVlTiNftVBJEVllV3NKeBRfU6JIq/5GY6sEIE7WwY/t6x7Lkx
yUbHK7EEUD7HcBaCZlx3sO3+BXMrLjHpPa2UOtyp0WiQhkVGTuYhQWskI+FGnm7baKlVWA5nnQt7
Pb1LHLFsGVzNCI1I83Pdd+4G6q808jWr6S8WF4LAWR0MdIvkjceEtEDYaCNJbM5YZrVhHEmXxDWX
fo4ZYOeNh22AsYb8Iw8lXj0FNNa2Lrvyw3WeI7tQMKbG/n7RY93pQq4EEJV0nlxszQYV9TufahaB
DF/h+FcZUN5kn5CMdkAVDRQhpWlo4rGIPNqmk1+NJ2fIepj0f+g1LGGVaUNzDsAn3Y0GLiu6fPOu
3Rfo2dAYSdrPeEX8mpt1HXO4R7SmANXl1ybPzOefF4g7ZNCgervfWI49/Z+mkZl07e8ERQd6L1ri
HPtlnVBrURE1D0X81+xTgqFFpnrHjBcFklIAssW2MR130diwHBvlxS9uLej6X05FOLlw4sDBS1w4
9kn+Oq97xVAPaZOTDG1VuGpqfI/W8MjNDvUMVTHDUIWewL46wKntYAjQfTPEq2cNf89I48SmaLCB
b5dUB85FpViRuLQ9xqlpPcPS716SfVi+9nT9RBoWiTbb05B3aPolWYtBugoYcScmRjsRa15XLgEv
io1GnL2cfMsNPqsnJlXcJ45SecbMe/k3W7b2MoKkq1a+E1dNCsZbzZQdI2+daKVHalzWQ9aJ0SMG
GWCkmlY8qu/Pn1eOl1tejJbH6gWweC6eJcbmLf7nMcjlfjsvf5HuC+4t5JbnlHpiNpYbyDUfyfiR
gvxOSn4VIqruCeD38IfkbQ0SnsqAtxebWV5oREDVZhX/s8CsftFwIVZUqyRW4BU13liRhGJtFY2r
mcLSvujZXbVwwhHX3iPadoIV15J02ucFdQxAp7rzuHC16/g00mgu7YY5wZo3Hp4nSLzBhacnlDw2
12JHhBrcNcdghQ9u5sJGv65OqslZrfsY7CQjXjzJYcgCZXkiXAVETZ3/o4NebPR4/sCPgDyEh3M+
6KxSAzGYT8/hsGptd6iAZxxMIzCNroPWFcjyje9tazw6j9w4z3SlhwWWmN9onSf41ZgdIgV3k+d+
Q4v+x51kmHu/8x52mKAALcHxGaoLcPsbZ4bOblDVzqoJVB+qZaRwVFCbI9kiLax7z8Es1MNgrh+/
AFGv9PoELed3L9jbGgOGIQl9OweH4raA0dSKmulVkjdKTZIkRYqW3HxpjMN1NDoS21dycpDZrmSV
v8V2Fvaks+k1OglBw2njT3GD2MwstwSQmxDqlleqZOsYoNXGoq3TuoGur5FistPuKamxVJetZnpr
oQD3q5shd31UwKQibSn7II7PYd1nbmCbmP3yZq6bLayAkx09A6ygTEUdlC0wAsTCtq6Xyk6kRlPq
s9qYBNYpplVn3FYvztAG+e4JvIuraFjzVXU9LKHOkZsC+Iq/n6PJ7DJCpgp2PCpZmuzu00vzQYAk
0pR7q8LWEqrCGzuCM2Y2POpfUUzeEA/TkwSsEVPlekiTJ/VskXakePFv0x3YV8bmw1IkSCozXoIW
FmGVL8qC5eW4to9cHIWwxNRpr4h2mKy6cUZpf9NEvKSEghbBQxWEbdxk64nXSODBwOalMHDykSw/
XBJr5l0mYyfX/8qn0fA19R5OCPXGN+l8pouSqewq4AGrWLLpQhsJ8oGlAyahwgBZxDscFEKIRZku
u0CxzSNsdTbRViAsRTrotdufJi3aRnPR7Hd/RDFsEq6hbbD8q4aaX6yL+gvW0u4fC8z1B/wY7wEo
BdoPJU2s0a6c/XfdYF4ALaGLl5jPAUJ3wGqDphqhjGYHjt5cOrM09hKgJsPPMMVjSbDQDh8uS1di
9b5oPS4+4KHlzTe8FdOil7eXI4I9IvW1JQNb6wgYUrA7kuU4yZM0BrhnuocEJZfvpTYjXo1gBI6t
N6maKtN5oc4y0PHmlPgfo4PyrJjLYm83xIpqNUFPA23TPUlVugwrAM64nu+bA7yTiMQdsjjHIb/H
BIUVPMB3aL2VW1GiYrk/uhYB4ZgE21jLCQonUHvCJTp6OEMzcBOkaB2phlLesaAMTeBZdsPzgNIm
1m+xxcXLfuXw2GQY0G8PKVc733TyOnmaKV6rnex7/TrhX1AFnUc4nbYJvXfdDjXAYhO7Mc7zOG2c
RM9s7WP2o7yBysdkrGit82cXwq6F0rUiBgz0J3f3FDy65yrco7DYsgrIDGlXOzzB6G7KrcQGoa3c
+Ef16nZn5YuEXkctwJiW3DItLWN3Yqq1kF5lfC+Kf4ozmoCs1vepJtfExTgmxbiIfH0I42k51Sty
P9CDdBc+xjKmOoCqA6Af8nyBX6lsA1hUnQ9iISWay9cxxsyXy+xHhnaKPYz9YjXrqq42868WpJRf
GtQKTF+tLKvN1Tvhj1HAJZ4dqPHdQUg+hR/d0sMoARPU1gdfAK7HzfHUERP1KpBbSMMxL2z9n1jS
oo8tNfqkR67xBpGWGmlFIwxBJFKkomMNYbFpBUfC3Mt1hyrVa9eQjCzWwwZlZglh34dg+l0vRA2Z
Ovo+dg1Ct/6hNJ8cw2GaA1Q6OlizR60mLQJiX4AhTd3zCS0f+4CVoMx7yDoujxnHt3yn04NBiFmP
dnI014l1OBFBZ+jYyqGTxtUGCQ1TLoLx7lNnOqKoFpzV3uazgdRgMPhFl9zg/zoxAgXYMjuZwyFQ
OgUqXhQBytKb4qTkBHG21oZ8Ob8TjDh88E45ReFyHxxPFxwQiSdwHRkyZb/7rBvYYN/f5yl9i7vj
Fxxrv3WKsu5c9sGsRfWpp44kLCIdtowSqTLnXseYoLlNOayFzloCCtXfGrhA+HjLfteUt+GKAiTc
FNvh1NmqThvSR0r8jxfdBZuOzg7EnUcNo4fWgZlMS3rBV1dAhXHrNU7s+eEjsQAa80Z9yPiVNRuU
HJC4EwDst1057OVO8zjTRuyyLQ7KboR51yWHhADydjnHDi0f0iHa8A3VHNP8wDXWlR4rxyBC3hKA
CEUfChklcAmh7MAP7ywc40yi3CKpnBclNtcRd3sQhpXKnQSonO/LHywOFs7MMiZvZPrUfNUFDbsE
VdIyeTMiwlTqQUxAted5H+fLhaLrLcBcflzAEABykxJ9G7qHCwulO/vthLuMnw5LfFTNWBoP6OY1
4MhpwFW874glut9nmJGa8zL/dwk+Llqj2A2xq/uR0SIKM9mkIAG3VwBCAUMuTnWQllJ5qsFu9+Hp
8pFoKnjsrHd48FUuT5N0EDU+6Wa5KrjoNQ5C6SbefdlXhVMX1RTqqZ0bgqKRQS7hHK+FoyNRrNq8
Cp9bowgdNq0O//IQH9pR14/NKHYZ2+uX9E9sM66jnfmk5OH80ot+YmhqEOwrv8dwSrhF77S/kg0W
9bwHbyVsRFIRs6m1scrPdsN7eivhNsSWtc69Y5OFUOidn9o+ImJy7vnfxil9n4fCa37J3n6B804p
NKOyBlVafAiWinZlm0ysZFJqG01C3QuvTC5xZxHCqOOmiiEWpW4D2XI+ooLZ4ZoXIU9JsRuThJNP
Q1XbgD0dq3F3jb+9Nx6rAvDM0mJPbRPiFai+63csVdEC3k9bAbHVx7I0WAYmWNhDmpoBE+P0E2KG
+0a4Comih0NF0rAqKIR4XZlBgInO66i5FuN22J5cXU3tZQ8PdYfxSvYW87dBYwfWI+9iRiGKjIGG
4OVapEjYRvnh7JDwSgyhZLdoa5zMS+Lktz9YNFoZjudnCfnKsAIil6dNGXTIEYBwADP9yGJp7/BE
3hbPspNpny3+2GEsKU9J20MhjtspqdNm9KPLH81xXU+WSInuKb4dCCMGLstzFkgSuPTKoyTqr6l2
iKjh0KdUOBN0CM5C5ROLlr93if40pDy2jHv4W9nZx1CNlK/dXME+aPcth+xyNRxD/NAIyE1JnLpm
Vz2NMlhUqxZpLYBd0H8JXPsju6mfH+j9MCrqHovd9C/zxwYk44NuZT8Xz8kTZfOfBxzG+hQg499g
ZGfPjRvpcIusEwHaeB9zcxwcs1chd1+941UrNgyVqV3mp0ci33c1tuL/e4ypzVVqyRWHJNXMPg/W
C4CJ8p1ktpBUULZH9SAwEc7v3b2KAfu5XwCiDSKacr2PT3WQJ0fwXDJNGcgy6os/+jwz5YY6NJYK
yL/Gy+ykzTNJxTPWnihp1eayvpcR2BuFI2oFh/XGxK+ifns2zQScheYvNFVHtG51L4PLuFPzW1Qc
pw1yt0iXrjhE24M37+yA3ZDJ9GyRVc78hxHMwM6VQ+fV6eolatyZKmggoFzicGL8vAVW6HRMKww5
ZiTwNn9vQPHFO3byKejxRMx0GjM6seqXJPhPVp0eSg6NNG/JuG7TXlJ91QsfELzRubd27IXV9TTL
SwJ0zclgDG8H8SdZj/UnjLQYyzE+az8a91ixJaZHXui5M8AT6/qbI2v7GAw4UcMq++IiJ9ljnLbv
MUwC81I5uDO1gXpZVlcx8Qs4movY0/tQiJHfRD8VxGVSp28LTCtvIsRvrHdOOrL4AKq1ikTvu1Ue
GzeC7O41ROWrwINXGlfYgiki7p+UXoIZrhtA2d8a83RTIXH/S5lWtO224aYIWxatxCetK/DZnbpx
/N6zcM/G7uZTuPpViSjoQ6U9Z5ULsJ3pyxlVpyX02XR45RxXpio6eruEe3tjFn1vLhB/z6PM5xrw
RnDq4JRthkEmFoJdZ2w0fD6UlV8NErtIVQFERo48QO2Rcja9y/5ZGjHT4rvTW+OluhqihwDULr4p
Ky9chQCx7eE9p5lyElDbbm8wyPpyTPnEGdwHJD5nJNJhDU7KFool8Phe+4oBim67n2RJ+TFAmlVf
LbSForKKY+YsYcontpNZlHilBej3+DUeUbZzCfq03+L+XdgMWHh1dNrUYrEtTfa6LL9sBpg287Xa
HW5DCUFSCB6FY22hmkMBi+EjpkCyp4APjiGYTsCvRJ+imVl9bt8odrzsciEwaYDHjQWVQM/eEZmP
1EDpzbCXAQzZLXdqkIYOxyonfDZTTAsWC1XpJkW4NtyWoVFNlaFWbPKNenixwP9JmuyWy6BTBZHf
JvfUmahBMo1yLKkCiKb8wduNku338NR2H5cCFm8C5UH03fRDieMzcK5fokurFMmhW7EfYsW4M8+9
yrkGVpsvkaYvH9cfohBNrhqwYOx9L9o3/S91ZIqJwCqUSs38VGM/ArsGhJM4UIgi5RepfP5sIG1/
zV1jmC80B0nBRtNilk9nqlkiDxyGWyZpJR/bTeacbVMt5zdL4RRZjSBNBq8ABLmCJKxfP2sVjpZd
VidfZYPKzgZaY3VdwOX3po8QviKOYnCzjS+0h+HaqpVOEDpkF6A8ANutlFqhUV3lq8juHyCuORch
8jVNoV2PLWhZvkWwaojgswu3yZ98meJ8Jjf2M7JWe4L+a7Ia28LC0Xl+0JlL+meQPLfggVzQOnUB
ykC1r6W2SoLDpV5Mx0qAIDPSn5HkxySonxdeiPCE87LpggeLdtocRYS2ctFnZ4ivHbMuxS7z5oNS
mjLVR6mEfs7mdu/e6fXTHtiADY6SwGKmoittt4FW0oWCLLRO80mb++TlapeqxXD6EFVZvWHzirYQ
aLE8JAAutgXKKbbpKRCW85IvSaHQ1pqhcGxiEv0x1O7gpzPVpTnrM9MJ0fKEmirBhGTQdpLqsBZl
b/lXAag4YGwJBS+eEpSGI2hzAD6y4SLxvsjtkMiZ8GAPGmK+z17P905RRlAqL3qw21fRubBipoQg
qecuayJFTva2tPAGV0LBGMK/U1pxPwvZABZ0jGqCxDHyc9BpUC0KT6CXLFl1+5CtU9atnwoCBYuS
ZX+UDPJaRNUSUdEwBZb9h4VtaS68DTdmV0vQQUOmJQ7flrT1Z/UyEXLJGBTdt560/PxJumGpmc6R
N5cNfVjrPC8UXCHarPaZGvCKEb6Sj+Vn+yg6IIsj+HKumemaBuicFYAmNpiCDEQapyLSrsEC+kJm
dKTSDJykyzsMxLqjh8BOeJPo4p1DiIJNp1lG3rpBsAxKAB5G+8lVle3eBixUgnHdj9T4kIGC6sjJ
uNpb/GjoYip7yxquZLZjgFK93Gy5HzAJ2UcYf0OC8wjFBmmLLSXC1S9PK4ECthGQUW23w/sQ6g6v
a1u3KFCqQMT0dO5lSHUnagRM406H7c98BOL00Q0p0rcUTsg2amKuswQLUAGmshS19bN3NtYthdOu
gn1C1AB8gMn8XNmKCtk69S/oNPE7FQo3XaAoM+N4VRS+u4vE0uJr9h0Z5pk1wOT/jWVc2QRK7831
zEX4G3d8TnOgOzEZ/8+nj7ho7ovkab8vnMES5PBEsVF5SHycx4Zwoz09+RNRfKAuHRY/mZw76RgG
kV4R4HLpS95iM+tIq5Q/X6W+DtFrlu+9lqwGGq1FJZ2KY8kvIvlrmTbquv1NwNFa/vZtzoot1lIG
hla8/iMV/4RSW/DWhMPpWmyYU32w0T8M4ovJ5gAeAbCTIlBi7Byxp8JrVCpmBExwlvDYUfcljpon
VY+7+Gry9vZaH9j56XCehfXogK5IHhXdiXLgDM1PShnLbtug0Ir1AKou7rSoKV7P5Px7ePpd18MB
p4513FrPsBJX6McTfEyK3tMT80TMCGFMju2SUg6VWZiGuHIXkLKkoIp6OkIbjy5YoJn0ZV9zwJP2
1Cxws/ol60TWDfeoqyFWpnTfT2e3257/Z5X1usZQ7vv0kvOSyML5xQj7RQuuMqOkmpow8JxiuZD/
KPw3aNsjGdIc2T3EeAwc451fE05e3BduGcELsJnLXe8GqR/KmlHmuzhx/E5nmEWMkj5zUrYy5xj/
2b6bX3/p4DbP8p7gg0VZPpMygGfAt8r3qZRoYhKVc+jsUso5kszGF8S5qhbu+YVXyu7Ct6f506Tz
t6K/6y+vLcZWwu9rFxNlRewOQgmPMOpSovb/VNYD/UgdUQ55z5lmAYzJsAFy70LiR8oOCyODg7/z
K7VbFsZBPOwBRAMQPXezxxxVTXTmTWuSWR/QBGZ9Is1S3lf33Ug91nD3/pmOOuS/yHssn2sGypil
5T6ZJzhIlz+gSTxPrpqtn5WfRd7r21SdZZ0OzOrzK0sNL9ukGoCFyYtEV0yVeCcvAP7ROSz6kd8z
/qPrGImNP6DtdWYnEcBgRL338LygVDdmT2shGmbb4d/CIEbqUmEZveWcRwpvi5vKaCTObxAuc/ND
8pu0iU7bVxKnyj6A2EtP0DgnYf2qO54QVpJfhqYxRDDfulew2Ttrhd+RkjIEtHEave1EF7z06PGs
zxhK4WrqRIOfbK1p6VnULPOcoGEAltRN8fDz+pWLCdr8ibDfq/u0R9kJVohlraZS/aO4vw6cqh3B
N1IR6P3Js5/tZ+D+Ek+Q8JvkZg3sI6Okxdjf0vswdP1+97Hevbi1hKDxYMY054/CbMf+ir26mLHK
02e8T2ckDkzW+/QOm5U606/RgFvyNu0gPthC+wcdLDTCoLBvn562KLPO6hbKpgrdCZ8uluNGeso1
7ZNaGRD3QvI2Gn8z1IB+El6N+SpkJrsXJ/2ukeAJTd9cMujUAmO9le+wn2oXVp94ucn9/yAiCklq
eq/oIpAJ8ZI8Pex5AgGGM5Q5RZTxtDYE7qROkfNsCjy3cPOLgSPq7h59+Bb8Oe4x9A7lYuR/pFQu
O8PaUBpJPGptzJcmm6YHeyHRbEEuGX4QWcjp1svZa8iYKsaMy3FX9dkXOkNfh1AaQYciB5S6LA/a
adfTJVGL3rTNAfCFY36cPbYpIWXye5R95u9scGADv2rH+ysC3HA+XZ4mo3u1gWsUJEIHVNC9fU7a
75Ols1vHRsvQO6YG+H05OrvlqzeEMTvGiPHr4283n3UILb6G9gtUy1vxYRzVuQzQftszDEREPx2U
uEbvtgyZBSIwCaMqyMGukElFyATrFtfF/WJtIrSaSI/GCBpeB89rBA7I0IgP7WlZSrb+3eeEauAR
B9U+yWVDE1Jb7wZbynhvqPlr6Z6557nJ6Wz8VIq/Up5SsHeBRFjU3vwcyrdXDLsq3fi9AorXuyem
/QYQUZr8018YAed1qn5voU0f3lQQSjGWR7M1wMUclHiy3FcwRwqX/0R6dzNuFwK1OEUiZeFFEmOY
l8eY8gpwtG2/96oUk8vrOCMiYX+kw3xTgJpg4walOfYKPT6d8wH/5mavUIe98KCLZQ8s86WX0aMY
K3aYPjiR39IKErHh49yGdYolzwHs84xtCKQE2xGKMfaS8w1xsn+zW+ZBEkd+jg4Emu6ak9UwYeAz
AzaYQwBNRBPlZ0JY7prDIEhKy/afRk2qxIMBsM9KcC/50ESZ7+TX/BZDF76wlhTVI8PYG8OlX1Ph
41ePfwk9/Mr7A/HQJ2aa6xDhSp3bEoS4HAomCK6sknNs2p12ZGmEOd1twQ8OlbRaNum3oYx6NLm9
Ojk9Xog/gByIGCQGIgnRkkjwlnpvT8exqDdRNEsk2FOCckqwIM1bGud3kET0pSKWrXGQf21OOwH+
zOgKXN9DyobYqsA1KCyN5C3Mj/6GJoNxVHtoteXlTmPXhqc7sPevLFcAwp1B0LYc7AHmB1GiWNpp
iMmnK59MVErsf8ab1YnnQJlSPEtvDj5KQLKFG9WZXnDPBdbycxOS7vppeaBeFPEAZWtpOtKNg/57
/DZ8HjqCOlaG5GS5/poF3+oG+T8de8ylaKTxtE+yxiZGGkKsC1ysClzHXC9Wit71YleIp5d9kIiH
mw96s7lX2e/3Ah5wMoxn3xpGyfHCXsJp4UnFmYVO3e40VNkxvafFcYg9ob/IZAI/0wCs96BW1342
3Ftg/6IxZdFfHj2a9cDDkqyi6UL0mqaXoKbpwDDI9anG4+eTpNTi3YMIa1ByCxJYf4yRavZJ2QB7
rAxl9tVibd/YKWdhCsMeXkEBZm/sqWEmTbRwgIirQGhvwehtpnzat4Ks8bLZcSKZdKYtq9v2ByB8
mFRvXAWcn74MuQl4RxwU2NAAvLETrZtbwh+hbr8np0iSGMekB7VCn22NCxEvtJCYLcqwALNjZULo
7Am18BvgH6kK0ZKYgEGha+j17oIbghPdHWFcSmLNsy+YUX+TGl+1EcttZq4b9Am6BFegdZCaSPuq
4tPs3cKgpJ9BmU/2MME3WUb52I1fjUl0kNzMril89X9eKG0wCe9dweuthTZT4He1aC4OiGLz7TBV
TRDRJ3Dy/Wq8xzjUA2FLzaiJvhvkUfFnk5bMAnNEmOfuEn1RKaDXaHkWv51BZFPl9xHf3QU6mu5D
UlT4GDI8uNU/WLfG0oFGAEjpobViNOaBjA3Jf37hmoK2I+Rbpo11HLYiER/lwXCZjLq4O8HMQkAx
nSLoJoBciPBroFRijafQ0W+W41HtP6gzOwLKlIjTvITbOC+zIAS2IZjziBbPFMtv6EQoYO19Meyo
42aTz8fEmTqByI61TXNUZMatAyPDpDqx9KdD8aIEaT3IA5rOMjAqywlQot11k7Ou4AtTjuq8aYt7
tlWHEZFg8NvpmdjUwaLaLb954yWDsT7ZyYwsIc4Ri332hqoEvoAB++roFnrJU0EPXJJIGaOzcqXL
eqtaBZfm7tsOVrMXavTvvAaH62p7KhGLnRUBpmRre2UL1xeJ8aJdQR9y7i7Ie26NOkfrFS3NtvpV
PzIB74yVGKyjzfLTmQqmF5R+JwcVDMy7Dnr4zm4H2LOICF6l2t1PnZhGuCbrI/wwzbxWqZpX1gtt
+/oXoO5zKwNtozYhZpJGiT52azyrh/5ycPC4jCXevinarMBjRV8V28DokSOYeu4gsWNcIek+LQdR
X2hSHMrdGucgwo11XQz7jwQjMw71redmGFu8HLxHN5sHNYSEFGqRgfmi1cY1IoGdLi++qf7DtDor
k4TDXZRNvene6HxvcB/FsI+XF4KOp9JPTbqm2sybQzn9MnM6whSmrdvMeTInxPOHlEWYU2hhAmMD
hAX6VctNbZUbd1/f/Y0HCvWF/cbWKmj7IYUuX7MZHJ1neLd8Z6QRkCDcAJBc2dmE+VkDdhKwyKEG
9tImGlaXvF0nhEIYqXk6U+76ZX7UDQCdKkdl9gW8ztTMrjzSgYVb+r5+Xy05EB4E8rKsONwJ29jc
mZUfunyqyojyrJJQJ4aZIddRtWCTKCU8/mjz1AuqlkgHydpTqHyeV4mO/2TzmAfPcCYgFUVqjh8y
hSmEGxP5vvhX/s2uChR5JxUQTUulV1KiKeYppa8+4vKodadwyZmKJWnP5ul7WZpjJgeiKwYH+xkm
2DglRspic6MGqt9vw48D81DE6PArsQoijD4goa1MXOx9uJ2QIS6Sp0hH5+/iu0RIWxO7SpdzOHG+
uj5rRPu26BHam117vtmP4+8ZIJDdfjRdCeZiaibX1M0X+Fr5Yt6tgEL/B+FNHRAWPQPy1pmrtvfa
NzdRmICcXlZUfZuPcJC196WZGPnteslKzaKQSHYJuJYRixdr1ZdvpshlrQ4SPnIDq7bNWHmanjh1
IDapbTNS/6dINctwubEtfYnscKJ2f2QuKbuUpkR8+7Q5emcJIg817rdeol401mRNRNPuMe/GpqPK
+qpM6ocfG5p39DWVWoYEF0s2kzdpRXC0ZI9eVlcGCUdUGScCqYqbUKZQYWYF/WAQRu+7s4JX1poD
OGafWaIhvLcmeGNY6lwe4my2RkuVqgHJXSLt9bTemEzi8U33rzLoPZ6+nOmgK9eoZdIJp1clNsPV
QNu+do4yVTvwBTW8LrL7HmRAUynNerBIaQeOgS33zMNsws++1c4uGNUnuIzi++bt6OkeMP2QiK5I
SPISXt05aiXuk4tNka4NfsFxjfkN8RhMev/RmKfuu2cMdeR4jOOusiwufJ0hv0eMu/OJB8u5sSb6
q4y60pDbSU5C6te4x71fS0lFcI5C4UbJ+bKyvwYEWpcBsH3/3JmkJUwFDfc4cSnbkqY2wJCHI5mc
WSQXVXWoawUCE4xrdtLriA1H2FAUOQMP2B8dlgO64rQjtx31AAtWfxcLLmAuLyUUEa9DVUirA9GO
lCE3+Dq8ApEr0N4uM9JDNvZzkLPczwKjKUqDaSwj6utT6QPTjryrT9WOgUsOBYGN4TJx5FRKHpCM
qrM3+M8MoxjTZQHf6/S0ztA6sw9xvuanMO5WD/aGIBFKMOEH+8liZDJ1m7UiXjHV6pv6bJ0Dd9TS
R/9WsOLBbERLZFd7xRCLXVEjw1K5oonaH1Gw/pUdqcUFdZpSeYg6fR8nnO+ZlXq+rryTijJbW5y1
AlfTVmS7Acsw1MdxPRgz1qlRqOeC3YZcN32hzcvOP15gV818J50F0sBurOwwOvTzMXqiuerjaBKx
SCKfPFFjm2FYqEwwNgtM3PODeuQQ6WFQzHBbkpnN6BT7CyfywBa+08EFJBHgmxHBAkVvj4lMsH4S
YrP98lutjxj5LvtT1ehChqGYUtGjMfr9mX3fDsKdQ1Ziwj/0xKgxRwCsVW26soWV1smzpX/7z6y5
nka8bsMEprTx1KZ9i7DZecLYuIxUnAxaJjJpaZG+RPVtbiKb8yZ9n0oesdlpteOpNT106U4R+e0I
I/FZiIUYriWOVzkWl9huMcmpTp0gTsiwt0SpNOpf0kwDYn0F1fevf55zOIjYFAJl/8GO6RilcnoB
vADAYivrfaVSMV0Ga+Jr7OnJdD9iVFfX+rJ3SA9+9QcHAQ8LmdDCFVVAALE4BgVcta+fQ4dryI3t
lfxjl1W2hBIi3vA2xi2foua7n49XUm8jcDHVyXWJnN6E3X0A6z2CdEtsPa7VXQYF5pAx+vdyCdEp
PN05t5/xda7Nc1Y1GSLwLd8t2+ZB9EQh/JXRdiR+XE11htLSq1u+7Pf+8Ij6tTRZ5Rigv9W2qRdW
tY30HHbQ5Hfo6ByYBiqN+WcQb3btMk+jRWjIQ/D4lZxSQtspYnp+VmyLjCo8ot51bS0jzg7hDnPq
uok439xWI2wG01SJqXvoqOyVzqfmLe7d5Q43S3B//l20cebLz9U18+BmP2syEaGt4eghLJweVZhm
NT/x0wWqA2LA38tbY93bw9gIW/LJbd2yHbbj/e4RsrmMI8gb3RDwKk9SVd8/WgWolq1B52a+pF/n
TX49D7SmUjUYnTms9bVCe/xulFjC08lDuEwqZC/MKcYPiZQt4ZnTYN2BRtBQrMkuFDYBPRFLSwPT
NcBIte9UQ5cPV5Hi1HBlSK4+TzqkmeJF8y5R7BxRhPAgrM//MGMh6mG273PnRMmVNM8PpilVYDd3
tlBXwl4tWfhY4GYVsyEjQ8Tf9EwVh9JVWknfWdZ3emyL5HwgC3V7+dk3WEUS2ACjMq5bvSh9fy7T
1KH02BGgws+/fqOcN0Dx/wIBbXyVU7lLUF9WxYbtFN5+sGCf8Rtp3P27wG+pIC0R/w6gK5TZJkrG
2Uj1yHEE8vRjnL0xc+RMpJmsvqT6DfWIAvjcYRm1joTzBWiLeAiGIaTNNngaYqNbk+SMMHgnWjO/
v6f2vp0pzkOyFDXY100dMkF+2DtLbo8o33mgwWt5IY5XynSGbB3ERqFc/mzwd9agHMsvv251aXWO
aLRK3ndFJjl52h9IcbYatrv6ubF+n6CYSfc7prhJIf5dqbJ13Lf5bALmJ47Mdqc9ozFn6o8qJ2xN
fKtwJNBggHCKfEMkZXXCek94CsQUGy2gAutmQWgqbJbzOY+hjqridAeX/sHvpTDjYN7BXlFd1W5/
vVhegBjP7EMvrzAcEkW6hY0HNyksBr+8kAderxLnvwwh/HCcl2xXGu65kdBFm3r7VzD8au9Z5VDN
PFr67qcwCP6qhHUZ+uoMa6K5kF4tvBgqAPOGvjGg4BqtSczqbGh40dsrEbZCKcpqDvH8zQWRXwQ5
cysM2NXYIRSovyjmkWW8nR/G6UOSn8ciuPpZKvLTHl5gh3YxGI5z6fMEV/O4kOVyCddNwBal/BGQ
H5GZr3P3p+O7PuxSyk5pgvOU9fkukqyWTZC6oNq977SMD4GmSfOpOFVGypog2y4xS6srrkAGWLyx
8PXZk9Rz8cOopjn4u35Yvhdj0gXZ1fjtyA3alpu7rG8xifHaoeL8gRuV90gGKe6hH6LKyWyOFjJ+
MytNyyg1OTpckenn94CEyK2nVW9imVaGjW0N26GEkMECy9uRhjWdofeWKE9IXRmtbBgnVRJWXFtC
FzkVd7r6Zab6agMz0f7lB5RuXi9aQO3CWv8y4VYtW2TlCFVTXxXsgBVb5aOTs8k2MPNJWvJIxz0W
OKAtOeZCFVmatePYKfeEv8EWeeS6+ceyJf9sKbR1ww2oLoWd2PvBZ3CJP3dV47sdeH1uFZ+M5hpE
ZtGTvvfOe+0/W7R3R5ryhvKFh8s62qWx/ZC6i1+wU2s03JFGd5jEZ/X6KNWBir8naVp6yjwrpSvs
AqzQHK24IKMyqux1AM0TszOwqGI7mPvpz7htslwM8fJjBz8Uh//YLWv6z1uI0i13tYkLtU7ajXhC
MD3uv+iXbo+Ty5Wj7ZVLIJ/hHS4i+QrnUZuGradHa5UDibaI2MhAoJAoTTezbb3Yjn/wYkO4a9+p
6WuF4a6+Z+BhQO0gMG6DLjIQslS+xFdOTfp7SDU7Arg5RNgnrNqlk/hAecng87uS1URg9n5Txim0
2ZpeO+HmGhObgKSJ/MaMVUvTc+RdobWmJNNrw3f7xGaXbf2kB49NogxXaPgUeb5lKO4pS1Pq/Qsc
O1jFMKBL6omESDCi/NSycLLeczjg5J4I0nlTTyBimZMTWF4LS66uJpgfceojZ6LLvuKLkSuzrl9x
SnGsMVwLfcSxhPjXhLMX2GYfbe4+Wl27RsdKmpujHB6IwehncYBM2CZuq3IkIVr4C1ErW86PF6lJ
Qv0oT4WUlUh6jG9/laC9tbGc0fdozdv06SnYBz6qaw2hKLM9SD+av3zHuRJ8LcXXkdKHY1llJvXb
MBBgTqubMQLCMT8VkXWQMG0ftL8JUgQLp0ZJxMZ4jHYYp7kxVVKwTzfhJbVoaae0oBwdU1EschbS
3J8Nr/00MapEkTHln7vbZrBJs6w27nSajvcWm40MHa9eWt6G9B+WW1u1vgdfd+nTWFAJuIcb6pbF
CQriRFL0UN0FNo5y/YQQeH5rGhlMR4bPIEG0WY4fuuVWQJDa6iiY9igzdmHW+GsUU+KOPfN4oTgf
f7WCEnM6Le1pq1Veq17VkDw+4DkUDyG2+X02mVElB2bl59Akufdfo7pQvaLVRgSeL05dIryAHzGc
1U6Ih0dCocHWmhUtYVxzRyQgy58nTlI/gMd+3UF0Pi0KILgOiy6dt4tYW7lzFXQPy2NZtlnglGvj
Ukrvj8guc2463E5P7Z/nWk0fe3/b3oEyd6+DBOwjDpza5KnUFS+ojmSpB7f97cxkNTia/C352z5O
0Ivl+iMasWrtTTwzBm+NF1d/trpszjHs7RFYp40n9f/YLpoyLR8ally7DmDaTMH7qpxE5DeQPVFr
2ozr7cFt3IiqNIMQTuFpRZNnMSEVPGt9mZwBia59oU+WisQFivOuzW+ii9ayoNcirF8TgN1O3LCT
E1a8MPaFMgmYS1sHKsjLafXFY1f9REr1MSLFIEdJ+E61w7z3j3S2XW+1UsjgqYF6C8tVtKSVyMdz
/jOc9Buz5P6kioBlNBQ9pYu7ZLFTzbaolTnnBm6tpnPxt+ES6B3/hOLCl+j2LdNTqsj3fXZg/Whm
o1cvendLu/T0exjo+zPlpLV+PyAxRUo5l8Ozhu2pYhlkWkcbTLgaBSovsiG0WDwCK4ukSJLQS1RX
tUMamQlqwtKWZ6nR+FYJva13G5IkEaRACRleW/o0W4MM5yKs0jeqH/ZoFZDWZoyYy6UT0zJbLzA8
HLAqbuflQstjr2wdTuAePEr29zJetiNZ8IhVyqg5V93Yu/So3zSuDimFCC9G3z9rE+TFpOzGRvAf
1e5R95GcTaIlaLtrSpv6gtSJUqTxfViiCdLgQzL55gaCyVEa4pTdpG7DVrvq/zd1mhqchXFdMOmx
L4s+KEdQJRSiHHMFdVa4FZdt2toMoaYEVAt5MygGSkWro4FURPMg8WxzM/iEpJXU44Go1B1omEc5
8SHzwGTiBJX129oRduFiYmGYfRXUCPLho72MFHMcBa9/wfNGYd952+LQF4XTJ4ePwBbmcan+ZiNR
bQ9I56BAqqvlcP8L6icPsnhwE8XR1Fbk1gJUkaxo5H74Kr4jGDLd4K0FheQehVMbDMtg+v59RJMc
0XGu3U38Pph8nZZQXC+1qZGP3UMPhjk7SKGMkk1L8hSTRITQ1SB7DZP0D5aclRDZuFv3bFXsTHpP
oyGJLvEZ1kBHd5UkNKOnl/mSyoLOObRPxMGa53teLK0rL9Q7Q9J99EvrwEU/sSioH8xErgcOeqX0
HgPJtHQRW8kPJL8sB0ol4L9xSYYpH/DL8t8NQdSdEMD4ODZ1tkVf5yYZhPglg348i7Spm5t0uZZL
sHy2m65qsjNXt/+Nf6hVpRcsmRa+bDGvcwdWL26mflSFVYHsdoTKLKWnKwelurW+J1vmcyyT84mC
hd2EwfM61qBTWvEEYwHARR3wk3vf+rm5IWxD1qRKenSjc5mxuORPE6Rpi8K/5lJhA6xkTeOMD1Gz
EcKXxmBWxj92Xdetd7dnc3cNlxcrMRssP4PfNx106Gumgzsa4ESYGjPfWuhjlyGxKTUXR2Hf02JE
Qp+U/+Z8xsFCzp7cphGyDS+j/igy1drgUkRqixFdGKjKt8uT2jrt6wE++XY1O54myYN7YG2Kitom
/I60aRM9+xVb62R83BuKnu6GnkIhCrht5z97Fg4YjGPzHhxt3PT9kYbYwNXIQ1xPoYODjNsDk2f+
Llwr0NVAOUbvQDEVZuIDfvChtowfzm7xIJ2K9QtPrQEYvbN4jLPFMTNOiL8hQSsLLrKkD2kqqQRJ
k/Y6aLACWNBZff3FKUej3OJwZ0V49fKmhVTzVaQ7SyGBWTN3c9N0xqoOSDMvXknUyV24SATV+J+y
TUXgybJSntXOmtM7++5Iv0Esl/fCuKstwr/o5MDJVkuA6H7Ztp334za1QMTH4pBDevyovR+1SBJo
EuGvRZ2rB86A7+dyKXSubU41hrWncfhneINfNGJPADaESwO/CqixjJ4oVjp9P47n+8MSsTrviVvw
9gabLx6nlnIxL90LJEzgDw/ANAtdwakdzDS1qrCMW961K2MtotnunKAcnSXByoPcOEWnRGCYhK3I
UoWLs1/ZnoOEzu+MEyvu5wOLx/mrEdGY0V9/DHX++4EO1b4rxj2bgEr1blsJnxr+7MGkDkwXFBCg
FPUPxvPbIhxxzSbOCi20v1AL8GZTmMcsE5AN740S0KbUFLy9/UuX/KAHCBcVFGgu7socfJ4K6kTi
2oE2MgdZij7lVeYlWZRfjOdo2lQowj/0sOFrWEhT94bvRhfAuK/e5cWI4m3ARDyIjLBEv0ASGy8y
Rny128rcZbknx4AN7FiBf14oKovV6tpMMcDt/HAcZPO+W/LqejJNd1+3BeRe8jx5PV5M9DDydxNf
GPF0thAwAIm096zUSyXOoIT7L2DI0fYv97frkIXv3J5JlZfie8yoSEkiNzL9FpUxrNs/qC62s+49
B50DJzJ/jKjp3DjtaUu/9JuIrUixlvp7P/GRoKOA6fbN+740HlknvRyEwEAjM8V5NTTaXdL6mHzt
3Z7wym4cXUx8qS/UTGE6q3s6byJvAyMzDbDftHGkOhZSgxsxdrifOOwkjNhyyZ6Us8qB/lQPkT+E
hB8zpk0qz0lSxWDCTtU6pXGPEptkcsNbGAkYnY3pciHHMyMVQ6TR/nwMuEckRXWjQQR5Rkr/EKnA
YXy1tQhH1GtE7Nz6Yb7mw4BPRODyHjvxtWcX+0PZJCRyobm9Vabc23FbCp7eDsAFkjyAYZj1+VcE
GQxjI+7r8HEmCd9IazNeqAPVFYw9NEDqGnB9OtzEXlR0G31h7iv09hwdDTUWzzwJeEx+pCHRGmkw
F/C8OsutjnW0FJRnvHcQG6kfiBjiwxaoLPMMvkkGu4z7HqV+cgl8VXWz/zJVZH17qSUk537H8YfG
W5TZhSi3U6lfKzKzqH9l8gxaNwGu55TcPoqf9L5ERTX1BwxcqRLDbfd5loKC6bGT7tQDYhdrNhwF
/F1N36iT5SYkoG2/yMe1GWHwcGk1+3nmaS+jS+UJVXYpU/Ie1ZGQA/w0MLbA4XOLSq5qfakf8LGp
O7dIV7DPQ/jJqTzzR6QmyByTinIEsJDeqprAlyaCgIjqqE2tXkM67v2GS6k1cFOJQRPeJ4zjYoKU
7vwn19s/0lr0DDxT7zOyJ8U/hFVarrpNgfKQb12hEkla6dsw/fT6n7WMUc8Nk2Zt34KLtQ11IH4E
QQ1FWmQOsgdeoSDlGBTAWQuPPYVVDTGtejV0SAtL4tFk4Qlg9b6g/4X53l3EIPsA9COhUwx0ys1U
DUEzl6OYra6j7F/UpIpcyEzhAlylx9kBS+pmb7cFKQhSE6ac2Fmqt64O1UHFSBEMNsDoQQj40U6J
8PwVs8TUqrIjfclo/NSureN5rIrVLv3jEfM5nS3GpfmxK8SSCq27a1KHUZGn7RZSsjDinC2OvMee
JC2Li7Rspfi2a0v982Sl4owwODdS4kNHBc+80hWvgNGxA408tA0edSJTDDgniPBmQ8TA6R2p2ZMa
NG/nkc5cg14m8+EVObJw9kth0T/Kd0zOuU3ogQTrlVDOxAVFZtnwf/OrnFwXgsgiB0RNEk8RWq0x
2Dok94NaCxbvcpCwyHLKZp8xnS3RXZjW4dzPB0IcbtjXSQA8IB5HAkTBBT/0xUTfj8eohJk95jDZ
e/36zCMlVocEKrLGl20iJpTc5hjTsQsBrPJD8fO5wZp3I6lsfMtpMzF9KVQPUTZd8fLQB/VEFurK
2YW1zBjPwhvTKC1iciapC3Vuff75EG269FjURoeR01qStr59Qc/VD6dz1q1rAu/ceRBB/XsB4Jnp
vBLES/6fndJn9PnHprro2AvbCHKqUgnVWBOgX1jNeYNKgVXX5ze4TTXkR6yswflnqOwbDSA1PByp
9zuf2/4TKoEk9J1o/1ebOYNEQRDCHb8vQRcJuDvnOm3nT19AZ40hVFYkzhy2kElE3iBPoPPdp5RV
ViCeU7DgYqfL6+yU+mrFIWNwK9yLQLWEBqBMmE0M9OlyZcVRjnViZDvzQ5+cp9oYidYEaVPfAlgr
exh6BhwDqQOJQHi1xK3/iU2Ua7YRiVW/DxnpnKfUHpxCD4PDpzQRPrwHSvCDAeM9Ethx6WPzhJkM
NAnGxDt2AOTNLz00fvnlbxS/wYm3ssELdWK7yv18oTFkgUty9fbwSub8LXXiB1FhAbi6yNw5zelT
SLI7O44f6Xo5UlJvvwynN1d2JSQFwDxLzP67FSOXSAQbOJYqr9g4no4ChP3QV5FA2QtLtR7xsnT7
K/ffgHI8CC9PVru4sCT7+IFv6QgQKNt4MARWloAD+KJ3bqA+ueOQCf2GFZ3SXjZZw0Xrlxm73pct
v8lJdcoXl7TXAc9isnJUmKStBYTuDvFB8WFfmLHoqDR1bT0P84lRnngI3kNyi5lt9OHaY6Nj9t5j
vQVlZCuiTBUq5iuc6WvJdZtI6cX6PImO8iv+BRrDe446DSUDwcc+wgQDDpZDJ4NGpsZSyS8D5Vlq
cb8lnLXWUQw0PINvAe9lQt9Q8RMRHL2+q2Mj/V0xywYKoK1TPelyiF9Fy9JxO7F6luwLnGhLlLQw
JWFNbjfXg3Ko1TC/w7bOybktbPBgPBBd/6M3zgKqfojep2OkjvHk9qWEir5WsKuEu2vR71HwCPoE
3JDpZkw8itBTVTpJ3mt5jAfjDav8pRoBbLa/hnYS8IRkRPETlfSCR1j3grN6Q69x239EfEzznkfC
TchfJk3oCKE0ftvM9BJaubZJhEQxy3RYVjKJZknPecflnnxxut3ikuDrK8Ow6oyvYf04WISA+Anw
0Jf0XYWT5XolA/FUh+JsHlpLr5GnYmZdjA8q7C7Ci2IgC7oIPVwZUVe50fLz8N1RtoO5nbgT5U8p
Oqwp8Dy670F2u9S39Nq0zx9fuImtelcu/u+8nUBQq7Mo67GrZX9UyHlL3j9CKk1OvOlp6Yb/ZJla
8H0y1E1jmZFe0YG+3lj8LhqXjq7G5iIw4MS7DV1EHTM/6pcOPQU9AmVc8AjE3jsaVBobzHeTwhvt
WI2B585mpvwO2N8TWKrc3CpBC4P5BXQav3jIlqn37pKKZCNyJ3BULacDYelVBKmyzD591R3u8yrU
3jLuuDGcvyNP0u5Tyn8hQrd5N47MF6JVzvONizA4esGJtUMCFFbFFIswibIwn4dWtmZ6w3pANwTI
/4QwQp5dFEqUiWXlzGxgjg3SJh7nofJ6dZegNsh8GW3OMgYqoHK6W8rZHJeQYJRedi+2jLaGYbfV
3rIAw5CWQhtVhDYTdpfZJCClSi94IfDFOG/80E0PFbdLx2piChC7LSljGe/iwaNIbA8w8+WN+ugG
vuTaiFnmKe7NSr+jBSePKP61Khf7pDOG7VF68QIjGAZaIPrey92yLmrKjiiiW37ej5G3H/HZCGIw
RpE5whPq10lt3cBMFWdv0PJJD8LcPhQ3RYO7vhgWxu3naV4FAERbjMylwk4sD0wqc8seTRhriZSb
AqoevVXNdMZLi8vSw1zZIhh5o6ZPiqrscPSL5XEFoJ5t0Afslq2CSyEfDaTJ/CcNMJ26Gqa4IgVf
kbJ2Vn6i+wpVNpQgRmFFldEKUFh8aCbfaNWdUFTQz+dbimFEggE7vCzGwvrYkt1d+LyPAHAhMbFI
jFinj7rxQI+wiQ0OdtY/Df+RMYO+unXD/LITeJECT1ktDuodiZqQreS80mzdfVMeP47N0bzRu9RZ
tDP6AOs6ojQeeAJ4BnEuvkWUYoXnfimr0d5s6ANn6LSDRJTUp8aIQsg/q/P+yfeWX56bDXguO0L2
xFENT4QHvRwUG7/Mf+L1AygLifazlGRbKe5aJKTwbtCCytbWhVPNMG+NXAjw4ISAtLtXjThf8cLg
7aU+HvFtwUN25X4I3pfc/ny/DLsjctVfqOtPeTtKH2iDMFRZxIQwCI46Y6A1yvXttAK6E6FwMZia
uHnTcOY5TMVxATSiy8uw4TNjkEC6DtGLTwkWBvuphDXv/GeXgmIpFPADjnjsG2uZSALlzz/F9D9w
0cIdkZNian9j5NGM5GCLRO74XXwnBmXtY4d2qK3gUMp5l59wmndVzgKYPwpBxYra/Oo2h+hdaYis
7tAvoFA7H/tlwsna5DVCEw0A8xywAkNjKUfMwG+GMXIX/qGMzKVXq7XgORc26+VMCyDmVBJGiNL2
+DW+97A/de3ihYHpG5YrWx3zDkk0J2awqktZLc8Osa8x/6m4Y15K75ktFVhwUV3xVB2XvArtps13
VPM0lPYYotQM+6AqHq7+iUNoX8DBz0h5xpKXoifkvdT3l/x+RAc6e4Sta0JRWCTQGIrqd+iWU/86
0oxW6wk95Lcc7thRil8uUPGN314MIx4o7sMOhxKjLvHPNw3PgyU1wWgaOsRo8G7KS7HwYNmNuz0X
h0hygDIY0w8ObVJD9syFle7F0okYNKA380kdD8pdY42jE4L53x4iDYtW8g8ptXeNkBYaH8nxY2Qk
S0ZxSHSbwMkeUNq6901hq9WD81rvFwYT8sBPt+yukCR1AUhQCrNSMCVGcg7rkx8tnHftHKE2/5q0
kXUybqGoe5uUgW1CZuZaTUQ/jHqOx6Brr4qtFn854epT6lcWtddtOPnsGdyLcvEUC+wn9Rxkq7rW
FAYiUI/p3Uzfh0eIqd8kJbgebXL2Jl8QGmGAMnGQuUZbYPs8fmzXKcL6qa9Lx+M2iRBcGhdqPj1A
VS4IH+FbeZGPkJFRwWLOzObDrFyHIqz1BGa2Fb4ExTqIgQgqPDjcER0UM/oT4KpVATfEpq8HApDH
YQXNqp6k+tE6ZcDFHiOnlFRT/7Y8+e5kFPo1i9KMdm4Rtzr9krVSVVQ+GXe4CMGdQxj5ABXcr979
U8xmffrBMU7BQxAGiUcZ5aA4E3Bqd6ukIn/N0S5yTVckMd0MG/Z6pbzVZ12OxCTQDlT55K2tT1VT
ciT1RdIjFrDdSJMZb8n/pC2l+XWPqM66+sz3BeAwQCvv6Jp7ezWHCvi86kk36iTTESYQNm00170I
eqx0juRqID1Vii4iV6ld5ZiL+pGb0YoqTHhElVl8ael35yHHKFWfCzhqAJnI1j1dZA25rqAQp3es
n4g8MfoYcHqfbeDJ70AJqobeihkITCx+OXedR+ZUxeIzwErjwoLoygYEIYD2/2Em5eAkcFI4F/FR
p7O4LWBPvAcKl/O/VR3m/uUbLmteeneXRUTN8fSUSvSim72XhkPdYsMrxuy/hB4cMKYtfskxPnLu
60j941pObX8snGT4E6u/hE3/phWrPuuOM2Hu26AHs7oUgIsesUGHph2Vw3yCqRyGYi6XqP22xPe6
BwLLCReZJgNmjE5dvIV8nbbP2hsWeOtn7Nc3U+Qsr47bqCmLW7toH+wCTdgt5Af7/0eZ1W8C94xJ
vsbMjw+3zEYrCYl2r2HWE+CapRy0bZg01m+DN+POjtD67PFNFQWaggVbgTsBx/Ck9Gn+E56mMGKh
pc0ZghbvEqoHL9w4xRAul84bqHEJZAJ44DZJIidIpGIlPcc779OxBj3FJmQ59o5S4NrXVfv/GgbP
fAUxE/RdSO1jqWDkOtOHg7YU5f15/KLURu1dLZHdAuCNHopkKsqi4ZKmqVAYuyQfoe3dHJAkHBJa
afFQnhCoXJBPt8Z2t6ilh8vQCrRwmvV9Wf0stT9tNXc+3SmZpmi57Csb7Txeo0YBEeTscVYqYdIV
Vr8XtOqPD4C1Grci1QCFehTXMvD3NxYo6zI0Epcnjmgl7Jx82rJrhJqBoFYLJjZx3+RlAr2EaQsI
PXayaHfGB7Dr8A8yaYoOgif3LpX41ESS7PolpNnUCvwQwQbNhR8GnKAKUV/YYzJ1n9fJVhc6bJWU
eKr+n3uXuQHXyVYE9HwVYPWLXxamw+wYV1OXkWemR9Db87i9l9QVUhqXBScifsRRuJTz1wQYffkA
6/D0BDmiA7BPS5dpAIzsQOdf8zY/Bbi0JkaWZZymvCqjQFF0iTyPu74ZnNsEjHtMwfkIaYEE0U9t
uHwz6w6/l0Dc+tAxLaXIt/Yo3DEpjvFyA2+A+eRUXGrr70CBCrxwZl70ZZMM7OetAmsqyvwpji04
4sLhdL3pL0ygv/eFMAwAGlTyuKNNlf7MK6BzZqSGLfLxfFPaafN3hG/1a3qqfHLQi7+LAkU2+ujF
hKWYIUSaTOpC5H6mCqae4nU27qg6mOOoGcMnOu7V02YE1i6ebypXnh2n6PnGz5YMpzSic8yeq8Z9
L999IxpE/rTl1qcuOnz9FTPkV9FKebocKR9yGjKWJXlziySKf6bEVDKLeSbTKSMbWSIZOFEJkcEm
B08ZhtgYPGczrGjQLmCmK9qr3FjQS2QVGN2tRqtb1BZTyBxuPCPCMk+YNaxEuCcVPh9r+9bVwCgk
EpIqHkgy4oOu/vEfr4PaX+4qI0yU+0dclbdgFFTASDur7Eru40lEroAFAGqEmA7X+vADrunZi10o
PfyLzMj/+6GeOXR8uJ//sstXO/MFTdy3xoTgugbR7wwUcT5vR2K6e2k0VXyjQYI11/UtZ3SgkPfj
xxstxy+KvhvOzYa+TgaOH5TH3viEF2lMAvr6UCLA6aGaRIHbo06iXdm4HLI1DUY83E4NgPV6NK1A
iRkiQoD7lN2w8bwvOarVZroE05zMMBPU5W4jknT13Tj4kIH4pJwWMK8hFtTN3UDOFYj7v6Wsesuk
pMKN7Lc/9fMHdLzSQlSZaj60dUIWraBBttobXI6LZy2Q8US+LLUN5XKotzpXh2+mpdBRb5Pk0a4p
x1ErtzTAdXH0c2xlJEklLgW3x9hd9iXXiwuxBZ6iMwUZTpN3EeFWoFkKFQ14C25bc4TmaBZvwjJJ
9XB/DHdXkruy44zFJeWnb5c3Eak7xZq3hgGQfYZqdsEVULq2KFEzEBWMxSabZCuRGfr1ly1AtXMd
aQ0eTpKiaKU2IQBPoG/Q2+jle9xuTD1csRv9LlHVxHYFfpxuOgb9l+lUIfbcjghiDtavU8AzAHLw
JAN9MhT77y5Y8tpUnWjmJOEGVmSjk/Cn9YUHh8JDo01NNdDpKqN1qLk38eRNFGri49N/sV2zSSWe
RTplLA0sZO+9eXLPBh8JnpMQuM+Dpuvw1hdsEojbEnWKnvrYIZMSvb65D7HvM25QWADTt+VmncCg
LlhvBu7WlRgIU2rZnyGBxNNR+IxJvsc1GMrFNpNe3OEcq3eYX9uGpRLp4REGlcfyfOnoypx1d4Yq
zcQrJ7qtvz4HUKt/6ft9xtKUbS9Ak+QXlDqRu9gt1MeY1M2CAYApx9FsTbjUCwhLSVmveobYndG0
dyMt0TChDEkHstL+dI7FNE485ZufPCqMi8rHBRdH/buprx5NpMXtyNMKffpba5XGzZcoNn3jI4XN
t7CHfryvD96xLq13cbYl3rBIckP34gsYMKK7cML6dNpYCTWjj4TBZmi0VkoSqKP1JdjaylydplX5
pOkNp1H4dYBHqaNJdKEwnhQOV0qB/O74gFQqdxic64BH196qvPJv6DbZgPCe5RpaGZVU6CoV605b
T+uH+awGdcAJlSzzPRvAgOx2SHyAExV9qp1xU7QGNXPMVqVS3HbCJb31AWLpynBtPFjkWMWcK9HE
wfBaMacpwkkG+PnQd2gEj6ZBFMPpt7cp2FPuL35fvAFUeetXhyvLuVcNGmbEfKmMJyOCe8gXpBuF
LnbaTdDWkg0uNnzfb1lLIyJHquYkgKWnAKrzIdh+IpLjyb7yxvYK7IQWIOcILC1ishTMhKGB2A08
teKlA933Fstj66UvocxtWpkMvMT4otz75rZKOO9LpQBiheOo/MJAHOVPGn3NlTCn7fpfq4ttSR/5
uRN+5/FfRg7jepiO8MwszsCWtzAsoHnAHF+BHwi70EaicfS1AOinl/lDH5EBY5pxCUbSE2JMxHDZ
shr+M5TF8vmzVqt2qTTqLliIc9vi5mcBOyhneawbo3yo6wVySGsucTxMoUkF4jeshwvKWYJbOV2h
ZudGuR21MIYq4HxlwkdPAbUQ0zoiPbBhEmWszDiuQIt7t0ffD9lejRS1R1a/QsMVKflbw4u35KhS
u4I6qqTvpYcmpU6GyAP0i72lLQMOFIOa7PH7B9R86oHze2ua2WbLL1gIG8txkLnMcBQlF/8ANmOI
3dLSZvHXMWkipl9PsR2fd8Grg+JCPLQ0rYnHOgEhaHxbV/Mc5ZlS/0Y5Rqk0QQe7+nNcvI4ulrBQ
zhnTmYb7yQ8wkGZOys4Rzt2DSyzFB48pcxY9UhXZC509g2BH38gYApvYmdFFZMiCrfJdxYYuIszI
yguxRvJkiZdGcyO4GLbnNRD7TjjjNvEs13XeYYanWZoCallASHK3lVPuahI2zH9IvFdZkWhasDLZ
a1sw9okjKC6pLjnb8IJFkWJyZWWOoQQLIHMo4VrxoVzmVDvYXZaf8+sCU6azzP+FcKKRGcZlcwU1
LXTUIsc39zOQLF9z548UCeCE/K1ofa8v+wUzGZYVFArn+9wMTNR3qmUW0LXyEmh5UiqB0Gu/6jJl
dNJmYzacrwqi0sfesomRiABweamVyaavZMXBsiy89tZgNVH3uo2T2tDCDCMzKmsierdbvdj4SdoT
FAMYTvS6gE6a5FN+iV04F9NM/ecw7M7zuk8y3KrpDWZovqu8Z104Mn3bZQk5UCuLHKeiRh4eK8SR
9uloBeWanvRyo1i+36RkKjYwjjTpwUlGHivSbxJZpPZGDorROFC3e7ZexPnQl6aQ02lVaXBwtbNP
YWZO2q3/AADrEvRR4a2qupJwCPcm71S/ENF3TaWxvZ8/aIwC+lIbtMVdPjHrpmVUpN8sAmV97W5P
Krda4TXBCEGxE+AZRDwJOdBXaLDDcnoXwk+oGiLEEhKIDH31HpDErc0nN0y1J607WK2s62fH+g/z
08UIvq9CRvkYWekrdH+018nTMpDj0Dasn6Fe+roTTFPLJ27gD094ZQMQ4ysNtPBtdYsU8cZ58qSC
EDA9eZkXRs3mOid8Os4bgPGRQHlluE34A0iAdpYIz3XCx4aul/ekiZ394DVog3fG+XbawqxoiL0M
A6dMuUBgapI6ritkUJJ5PtUPowJ5M8L0r5fjkmm23QxG87aCoD0u9zwJrbAwQnmutxjF0jPfvWwT
7Xrx8RcWHJxC9DZh5A27C6EiJz42JmheNbWYA2r5d+BfeHE6XokVPdTdX/667hMXu79GgdDJFMfk
TGr+Szn8W22GTBlS4Jv3+i2ACBkIPFc4t9mj5rMAdZuObffVX4GMLL83ZkXc73+/NEdhu2KelYr6
Igvk4KEYCr4vK6+4W3In+gHwEZ28QcAlQAODBCraylCdbjKz+dDKy8A147dpLzYp5t+jJqWBRSTt
ZEt41Kh5PcesHyGITjaXTdZ1Rng/7pksMgRKWiKzh0nDMwgp5NS/pz+7QrQiJgelXc+iNy7wQrm1
KG9iUUfX3e9j7YqbSgtyOqGXKyEDQKtmfktE0uyAUk8bACRaelIf/viUdZAefO7GFp0CC7SXJcNX
vBY7/TaFNkDvvRalaN/TRTSt9RpFuakwdkaSDh5Ju98Nd//86TC5RYwJomiGFdHP2/G1mLDHjrmj
UFaECMpoNzu9KOg6+uWo4ETGUfYHgiQe0tHorXcElwrs9bKs2MZqTtHvZ4gcKkmnvG3F4xY2ZIlk
jcFvsh0daNQquT/33aaMhj7bSHbcbgDuqDk29BmYzqwvVXQlILwatom/sWu5NZpIQYLIAIOs0PnQ
l1nsGj3ANWUkLs5kdblBZ1e+4hwdB8zoccazt5ZrhZ/dXcxoyEkdETQq8MKUGp1sjuloPLuIR8xH
3TbPv17YKpCHNjyLs5PDbJ97yRE6ySONCyN2dolrszZ5/ykKawFhYFEv5q8hL2Vidn4DTj888GRu
vt9tlgI9xI77Pptx5NnHM9CvK2NUfvczmUgdZaoNj3Yip7SOxLjKD5SvpRg6xJ6Hb7hGvcOqMFcL
rlvuyHJtslE+tkHw/AdZhU8Bg101OfCO/yb6uUPOHz+dogtOI0wfqjJXtknMepKHuYOk2wLUQ7Dz
M5CQddVqlUXmu0QUw2QF9i07wuNAdA5ZZ6TwkiY00c+DjkuSr79jRzZS8DQWJJOyCvmWI+NaCUPy
xED087VuJfR6rM7iG0dI+gMdY0wF3r0xqghWCqORfLHYIyNGqy50SrgeYayT1YbILQgaBPpWGYqu
bponOhMUB7nxIO9yZ79W+29wZ7P2gghlPDbtU906sH1f1i81WnZuMC9iy4Lfau189tSY2HQNpelJ
PzK+wSDdSuFOBuzoObY4VxIYxOcWHevG2dy8aD5x0lgxPWzxTXTrOX73s+FOm6oslp8Qc6xS3OEi
9HxJodv/OT8xStIe7whJ8nXnKQbpSFYg+3FOUmsRWNrbTRdFuVCN0Ka77iIFsh2mcLUtEUzLDR+7
d+j2zaovhmuJhP78thxg7hBhfw7TbaAsaza2dhDZ9mErMaj7bBGJmPRuCDEe4CntZtGA9klApg7z
7/ktRPH8XAQ/9I+fAa96QtpOuSbN+Xng1xsFTclTtOSshe5adMvgpvvykSm8iV5hlrtk1EJpCdRr
X7Q7GzSvzNj9ZKEfg8RqDqxWy+ayK0+7OfUdRDdr8KuXIM1KDUkoqudVBIvRekvaXtASWmnTn86q
9bVEal9C1CEO7MQe3GDlpeLT+47I02GwDzEYA5bJx390g+gx8WEhz3aiDplHU4ReDKBg9nyYcFsz
KjaDRCHPHq8oMDrpoLAn5s8z/cV4vvgBHF6bHNASXeIQ6KcFIX9djyKIbIqlsRpvlx9ITj60K3j2
c6ngS7jQ1MlU4M5iH1oh+X2c6NC8sTYJAt1MpBky02dhZF8DZOoA7dwOwr+f47NXubrfY1w3n4d9
fn1jlYN8BMURSNhxV47GHFM4Gp29hbAT5Y2IPJuVWF9Zo3DXsFALUp5SYl52MXBmefdl7vkETTjM
QUGrmvQ14ACWr26okdF3r/N4Rf3hVUNfEw9CjVaH8tYFy/f49VCE8fjtrElAU+N3YSJr0zmvnbgl
hzcoZtyGBKshcCW3E/tmX3XZDpsYEZ9JB0pzG3PgoqEI5NyCv4ZDT/AxSh+Mcf+tWDjOxPUyvskE
SI3BLQs+Xu5fi9m/QXCvxRwh6fvCsWTDD8Mc6S1K9pBPmQKt1S57icQ9LqxLr3ZWQybSAaycGsTR
zIaIGblLqpHiLgVGno93xe1XtjMWrSbf1RoDd6npr+Am12RtHSvqeD39SHSTQ9c56hRCsyJq+FkF
XFboEO9x/7etvjGNmRdxvrgI8N0P2LXxrvIvEbIws1Cz7P+TyzVSoh7Cwd1HgQAJHluW+Hs3cGzn
JOktJyxAlAMN6Xd7mGILZblcEq1Aipl7GwvS++KKB2VQw5x62KTqrQ0FgYqgO0CrDaAra9anD2kn
gVP/YVYGiJrauyKuoKZLxmZ9kcXg7PTwJmH6xihZikzWRCUyTWhmVnQbzTkCtxLZahiOf6ckpk/G
Hv0UTn/nR/kh6ITRiRQ4b64b3mWAs7N163Q4GlUL4tkEIvhK3uhkeRFvGUFts30wp6Y8Hu3/CEJd
yDhf8CU2ENi6Yja+Fp2mweyTUghIe0/1e0NMejioW2+RLU1cRmjc4vhpFaEl9bubLWDb7M5NLI4K
Y9IsKHysfxdIeQILfWciU7lpQ1+Q3QYZAaIJzYXiOTa2pb5dApbJKqKxLYkegpMFsfRMEHTYWgrm
EzkoqN6odFfg/g1PYisW0edL+mTyrALlDE47LZJA3XI5pUf1DNidXcb9+SNrh9CD5HJGv949XImH
KftIp6LLPpmPOHF6xeUFLSNKpRhuB8jWokbSaRUGePpW7bGhykCo9XyzZ2aCXHDvERNplsrRlym3
3edUocP0W/NEMHl2yiiebwnmRl8W5Ig/Jpbnx9WnBkNE10PXyzFKUsAy7laYIy7NvhrMJxnHjc/3
8/X+QfVJuOjP9JEQ/pTR/aOnqQ+a54xczgFDI9UpnZEZZYOoD+1ekGBraTY1o+8SY262IWJZyRG/
v9Vqm2tLJreXsJYsCOVGTWmewNwC2LZdnadfqSr8sNxadTr/n0inlqg13SjE1XMLC2FxmyY8pB92
3neOQL78fglBP7To2WUcuApy/lszW5O6Ulbx4kIBoR6NBasyFNELm+0sCCIB9xCqrAg4wlUBC6an
LrST0ROqRWeWVEYCy/NtEA00as6CIhP3HrnBaHusg41V4hOLWqdPay6b87z2GyR973j1MQ4Wok0z
PZu9ZMi68rI7iAx8B2zzmGcO7MCdruZSVrt4BFEZR214olJBSV2lzzkOkzKRpbUmbGVsLB4tMu7k
qzmXAjuESHRsVSxCUcV9gKIId+2ZvJlVChn/f79vhNCVsMg/qhb5Diltow8/K5KPq3DToDRmr43A
YunYorqeVzZzAUJV3lJy/OILqDenTaULFdtRzpdnVgvt0PvBrsaVCVYXVlSNqK1cVBp6F+sR7bzS
V9qZAI79O2mvRHNH2SQhAlkGB/OJfQXstU3gEt9wlAUxPzG8ARt3CIUIbsefdvH165JX6tGDnavp
RObFOoltlR2FegGKuUvy+27RyhHp0QHw+WaqIA7HvaXDTDbcRZEAT+k8XYaJqjyNkYq21+nqdJ7R
AIh+hof85DMiOOS33V5LxpM1qhCaEF9jWcFVKxb6HeX92OsIB4EDJO9gRGGn8lL6eoVd1NGiCzNv
UMgW6GyMG3SFDceyfK6rNBTQfnAywo/Di1IEsX7H41qH/t8wj8wkXLUO3wh1NXiFzLjxTpVY2MX5
zvyXKPEMulWQRKGYqivYaAPSoFLlcglQUAGch8C6QeZyMrZH2XuKpZ/fzJo5g83+j8j8jaide7zc
yB+r96P1Oc+9G5UKjBvFsFGqWZsGrnLKMW8nDZso3ZkMjnx/nTMG9mpC9NAEt53GSOhrKNSl82/f
QuOMVzHydUHTV7KsV1D2h5lKpgFykbCOIWWpa8SYcr5r7HB6xz9JDt4320IexJJ27OboPHAhr9ox
ziZY2yfSDSDcvQ0JdaEFp54dAG44z67tHOHH3fOKTVneBO+LK2Kadkd3Nwriz2I8W2Quk19SiD8/
zRNq5UK/HpaDq9ZnXTH/VV1lIeZ3443rHhJ/xzLXYm1ownSH5tpbhow0vNp07KAtE9PHvbG81hNL
mwjF2gBLeycvyCeNkjFEcgXu/8ZsqK4x67XQzQC5zYqaNsY+GhR3DflaNMV+cF4sVxRo1Aw/PokM
ZabGpNtH+4bQqf7QQVP5fdix6PViaVjTHVY8+ldBM02XjDOV4UI+fdPxE7vBU9xFGKsNr1BjTdcO
l3Z80bk3kTNzIawyncpE0VTu391KKk2g7DNC/kIQjKFUUbBELLTgcPK8yneZBbixudra32Ij0GbH
N+5D9q5V6pJBPHAvTsi1KpTRdkj+nGxTFK0qrItns4BVJbMdkB4jBAdi7cb8B4qKeu1GSSRyKJoW
dMz3WyKu0UIWt68vCEYRqLeR6Gpot411uDNNOAWnXcEEG4qA1Abvu3kiwu2J+Q68ZkoAvcji72io
74v9pGWsaL9M1CAiP5V1M6OiSLmd8gWaG7ejVO/hmNRFS9bETju57n0vLT7xbdpSBphsD1e9uHPa
8BDqhPlwZrxLHoqjDJvL8PIdYPfrcgTDmrICJdvOjtgzQjqRaTqUzd3+GKqa4tGBTMvOlPAvXt9h
1pN5l2csZ/OsKnN0dHBKct65gZyh1vVsD+6QrcI8M0qf6JuKFK+RusHFJ7KtkS90d5iWsLkNrCBs
6yB/n69NuSsCZnXXogGG4GbwuoHzaxa0UmqSONYUtMHnsYug79RqCdPhJrWYQzD4V4tT6W54nl0P
IorNXFKHQcveWjBs6RdgsV+J93K+IJSzUD0XllE6KqjVTEUZ/N8gmFgka1vS6hUGa7EJ9z6q5Ebe
cQ0QsZ2dHxgZO73o6MqzHKclqL9Dfsbkk2O1541C4+ZuVzfB0xyruT5pRxtCRmwf9dKRcdvkKO6j
KRfglWFFHa0wBIhyILISZXwYUbH7Dlm+NwLcjud5LRTVgIAE1U5ClEYtrQVj1xaJkjGO8KJV3rWq
y7b11E2Lo2h7qikd8fAnGKw2/05llCPyi/18m6TCifKVACjm55MTT6NxfbWab3Yw2uOm1HGFtTwr
JHiCl0KC8JUGph8KfJAkbT6OS3G2q0/+ylgIZcEsFcg1tzRXM6fLYXkeYi3do+a18qSh4V0Vxtb7
gSCfFWvrALu0CVh1tIJOvJ1rBes5NnM0dJgJXf8RQivSNhKOijC4zViAO/QWF+pn88J7GBtWB+Sv
Coa9yrRw7f3hLBHKO+UZCB5KITsHUuPTbx4s4DdgTQI1X55LHl2Vv3orNRyxfvUj2xoVT9ta9x+v
eTg/RjvOtIgAiz6Vimsv6kzCtknGEmL1xLmThWE0EM0vjUjiD3WeFr9OM0n3NDqX2REKrS7u1fyT
vYle6kV3dqBxiYK85/kf2TCjWvMHc53FMdhaBP41xa3ohSNaj8K1MJzuaobIdvuiwlcAukEgmVt0
mUS+hTurjIb4BZiQG9gM9t7tBI7stEqbwZTBJABYKJDR7cop7F0cY1xM6tknqo8nOgB58w2+KSiM
NCyvLFPZyCQfgEvEWdS9TVX9S3ni2SSxJjOGWDb3V6VToXHew4eblO3q7AWMj2ZTU9JQMoldxrvl
JnrdMaj5YnXST6ogXy0K+y5y834vyzslZvaHS+fGjYwZZdR5RIKaA/v47xtL+eDJzBQuqiLQc/16
QM653/p1+4RNOgHEwXsDJObDZZfr6TioK8nw8yEWQnFFUyzBY/HtaLELeKpBZIqIZ4hsY7SmffRs
ThYafJtvGgoMnIFHlG6cQmZln0HCtStzzvOpJO5xSp2+Q6dWMokU4cX53ZvjnDG6GmXoX1fhWSo9
0ysD7K2vp836FsSorayMkYAIf803nMbPTtHqmZjGDM7NZhluyiFm7hmilPPdvoyw7uGKn6/7bRlZ
Q+vxoFyWvBxpDf2EUDCIbdRsuYNkna3JkhAJq6TJU8yQgWldBlyA48bP06e9ZV3V3XMbX6UPdcLR
6BKDs+aWGskLDTVmhJEGEcsBknGrrlQ1ClpP1Fm7oNco8Zb0ih4DVz1MYs9KL3CTGdF21i5gqx/H
aIUliOPunxJCe0NroMPW/zRBgi+shSbF9aCKqUyTCn9ODya51Dh4/QhGly9I1WsALCf3gyG4MXOj
31/H1hXTqZc3eApYy0CnW1L82/IT1syfleBJwORkfWEkPlFr9e/5DNL4yJlSKelaZ57UJdOvsPtK
FBEV3ANJzsP9pYtGwjGAal4g2b0sHT1IYs9CPF3crMioqWw9/rKP8fK6qSuCcpucz6K7pV0W/uue
9/zgVRvLb1qzOvKyYHQGcbvs+jbu2LrHGPn+si6VEJDcsj29X8Z5sU7G5M2ECLFDTG+cqCSuTXKq
DViqhlCp+9B28lr9QOZOV/OkQc1BbEn4xdjTfU50ZbiHyIuzFfPAMuX1OVCegCSp1Ofk7gCVygX8
yRQmB7I4nycRgl8HSsUSOuGoxyPylNrEsUbylbdcnc7dlxvzs+1EXX1KgE87wNxAgHoR94O32BpO
057e0532KDsnE0/qIMd1wZufewgHN/UliYdwa26ZqZMw3ys+HG09uxCSlgDSM5ZJNklcbmMYjv6V
yW4AD9yIyyMEPK7aFYIC4AlQf9Jn4emq8/bbNkeMmbe85w63Ij5gjNggRQqCle9LG9FVa6NblCQm
PBklJ/rlqlOkfE8sRg0NTl+DEOJ6x/YUSSv4v6ei9HgC6D7DFP7jll87KrG15QFCO+t0CZKKE9Hh
6SlxfmaAEUzQVopjmoJFdZvb56utDQDpcwAnzW8MYRV24Nl8XoVARgLqPrdYrXRVlifLZ3WrFFy4
g3/lPlE5ujri/XasiekJtK+SQbUGdlu/JA4N18ari4CG0mrTq7d/+LvZxPyBlcc75DiGxSju2iaB
T8oewLJW3HPzZDIgVNgermLZRtedjp1D/yPDgW3NVWTNKnKuY8uyRRnWs5FjAarHZN6z5w4hRxgl
lMfDZoMIEqh20IryPkaWujSNnpeepX8Jv0gjDlNEZX3jruc/tuqq4AmnT8UFYR4Gh9TSgF2TdH3Y
+lNAnizujWF5ejsAKv/sns2E55u6rTKtMmth4xjpMjxonlJZBM677Yhg95OwEw6o/xvkUOv+DYnl
U3hmFu2RL39jYq87wcwoYvWdgZhf/2WvRLDPZTcZJucN64dmEqajGCXPsbHw4wa+bKYSm77O8rKA
gA9IRUOtjlK+ZNXCcLUvm9NR5FROJ2OJd6aYr3PnsS1h3qQm23PGLV6blMRuou0lKHUTGl5fjAkG
/HakJ/hbhofOBRMIFsjMTtQtKu1b58sKsF/wpaA95TQokxXhddGfq2+hEpePqyUkmUQNmsbw5A7U
cISHFI5lgo6V2uTckTUOQd/hB3MD/eI/8p9+/1iIfu2HX1wFYq+IusHTBwB+I+Xyl3O9F8iIxtzA
/flsn3PdTOXHCwzhe44yrGJl7veAHLuyN2gHUkjoh/zlo6JnjOf54G5a5VTbccjxHRditgat2zo2
847JOGVQyr7nl9X8miP7GUjWDXPrCn0avlMo1RY4t2EW7+RDRvqOmdcLmyyAwAk5hj+YmCPC/ziG
lWyreRdqAiao5IePx5SkXsa5lQLGqesQmDQjxlQMqhGsPchneq5iavsMZvsQ662JuASNyAXYy3DS
/WGghD7ReZRYtGDJqImzRZirglZ/LEDZAKFUQMWsh1nijbt7kh3EFXkWLLFXoFNFWTY8JFkPpKI2
1hvQ2iiFK5DF4Qe0vBzjX62nYZCQcl9vAJv/ffHeVgEP4LOtrRBNAjdLUVHB5o1KLogzWgSWZ5zb
l3uvJ9TV3UH9HlIJe5mIliC8gw8uzjn85GUsyOh5qbT++vPXbFsKcaePpoyATCmM0dXdT6mxSEAa
T4xlOrv8NRHpn9gNHFkpPfKD5kA69JIaUvxDQjpZUaTq+EAgJiqe2a8r1AiWxLrqhvGYBRNpYGKZ
f1IrWpgOQMOsPV2Op6zUVVTamqvBNgWmmRjXB5oRQaYh2F5ldbWLxIVe5GHhp5c/AwwzQ7GaGO+A
ngvNW5/hzx97BAppon4CCRYB/vG3FQWntcfHLKS1rj3v22pQPEVpUyZ9AtkgLCoee/L/bqczA+Zm
7lVfN22DYhkZ5ZGPcpM4P+ACnxQSHBXxpc/TShKYTsWNge3FJAuweHtI+tQkJsqLjWW48mK5Knda
oX71qNINaKWvPUal0zMLXB6R9BGziMJ0EIPBbXclCahdtnWfXrRTN6es0Si6cwS4JyFU+TpS3VSB
odGKaS4D81Cf9dXNDiFetR7e1576eI/6fAzsTXiB60MrD0Hx0ft8CR9Dxbqi6XQGmrJYCVptdmSs
yv2q/xzUVZyIOfh5RtIl0tceMgH5uerazEFSrXwoC4tJfM9aqjZRgq2AP5p4Vz2eM5YltS3PHUD5
YjjXc+buAIQGdm33qwP84eQ3Ao6Pa9qNAHqpM0/S8moKx5rQRmL8c1n0QX1Y1XxCkkaP/5Lt8u6H
LKi9uliveHxFjIgelvE9pUi5QT8yD6eY19cWsN3dFSOKO+OapGqCKx6h1JBSw82O2YvEUI8lIWM2
nTK4+d18h5mIV+boQEd0oONxHO5BVUN6X62SArTplEeYlbFdHkQ/CJTJaZUF+z4Vp+F3EmAP+rRq
WWtmjx6g54reKss89NaRlKZLQo6TY/PEmvcM/VEDcsEPZsXjTU3etlKbS9W05mXgNLEAP44cPTDB
lYWQ0+QN2nw00UkMoMhd6A+LWwUWj/M9kfPyn8+RqgNzwxBR/1tWiiBKfdCmbTEHrSFzykBvfHk+
5CUyNjcfHZOUNXOM2oAPjjWcx1WsfII/tmkVsFjqDABWfnrusCjrdh4ReGSBlWiqYY1a8BiG1frh
HL9ZUAioSWbIo1e1QHl9mmf41XdkNfHGI609k0eje3bSwFwjGn7bfHkVQjQe7dUXBm11gQrDUHVR
t95TG6lhj2NhwBTPZA+AXXRGZF9bFFm+TQJAhm4eBZkwsrk+xYL04BD+IPPUSXdF6EHCA9/QweyZ
8u9HxeaOnVhc3Y49ztdV2kHj6uTAFGQzYaTF6en16CcD7YVMs5HsQbhtVNNyF99EwBqA1ysvrcTK
e+H5WPfUOkRX9Kh/vMBXDX3ctVBGjMm04kwo/t6AU+P483INAAEbI75XeG9k6E70k3WdGTH21BHu
GTEDH30+z3ORZdwyD9pvjYDmwlEH8+R4ZG+IZkuJjgh041kz1kBQTfbj3atoXNVETGRBc3UUdDOl
VNJcNYZYgvatasCf0I/MtgOztMDU1VYO18ygUnIcrzncOAxLpBhGKnAATWhS7Xk4mXgJWg5YBOud
d/3ExEtedFr67Wh6ezLdMlGlW4Fd6WST9AU9w8zSeCAjQOrffh8SDLXel04O/Y3aT0LLGfi6xlnN
kru6qbzeGFtNBEAksljnD7HB6X0fXK1xxXz99flSvvX5El5MMVYXmPAlDaev9rps5nYUNNp3ogzB
rIkyD+wApGJUeO5SCi726cJ9ll9flTiqfjRKqZBFHGXe2UJr6u1UrefaxmWEOFamyDV2bs3YRF2z
HSdBV6aU1hDS6hCT54mKIfwc0/GYDmRvLfpjotgG9SnTZ/iSedEcKuE1pigm8EazR5HUHTbPPwJ+
LYBK0S9awcyDlsu1E3e24NtaOvbWySEqWSeFvKlcM9HBqieZNjzwVf0gD8w98KwLXmBwe73xwDnZ
3Q8VC2SyHTLNc5LJoTJbrFQLIQ/XZJFpwwCG6UZcFu1q317Tuea/7gMllC7cu/+4iy3tYtpNHXjM
jR0no4hArkLDxlDScB7XuvzUNmGQr4P8cDStzZfPHwKjwXaj2HJ97o3lkGhS2/FFcmjjT6hOfLrm
qhs/EXzu7Up+pQX4zhKVWdIPrjB0t0g6Wwy6RUYHhlc+tAc34FqbgSkNDhscCCqHo+0IJTPmHtJQ
Xt2vM4hwZJ6/Aas4F5n165GlND8youHPgx57lCVShZ6XUDegv+XiHnj1WNooyOzdsLBK3ZajJh6/
FLVTAm5uJ7HF/0crSHZHhWxvePBoXNjkXbXZr/wkMtyX3VTz8aq/ZS2yZJ0Br4AvMklA8l9B5BGt
EfaJznkuwDZ0F3hQHLuNSYRRbvKI5h/YknscexoBSd8qWLJYSB9SBm8PLBTove4reUwNtzd6QoYr
cLxjU171UecslFSMV5AhhhcbkQhSqDBsJyeTbj5LghlEqSM51L3hT4E+iIxAMh/Jg0fk92lP6+dy
fWY5mRWAjECFbXbHn423jt4Wym+uURVOIW0MwgJ6tC+dklE4oxY8rbEdKguoWiec38C4Fi4NfGgX
rp2GUf3/saGj9Ne31XjB521nvnAN9SGbjhOFKnyddwxPMJL6X04XQZODPWoua5gVisESdgSFTysX
P4NTTI1HLvLQOgNehrBPOTcm27EIDctMfKsr7f1L7N1F5JWyxa3/2JYxBoOTWSzjo89aPovn4PNl
Xjds8rLsX5tWWby/fGupG+UN35QtIA1z3yROIme+ZIZOTHdUYR8MvItZyslpaY2V1iq5jYzKq8uR
nKwHX94Q1UqiA4lfqiXLeQKE6x3LQFRrP6K8GXcg9tXVAnE1HWprY1BYWNicOoipo3IZDRkCRshM
GEE/BR9hXCF3dEjbJxQttPn/BuR8Js5aiCWn1P5KrmAuGJDAkcoJsxMe4FFHOm335Omhf4KdvHaj
DYQ+M6TJdYRlZoCpuNQRc/ape/kYq2S573bSIIyBs/JxrUmKCMQqUXW2oGS30u+GEBZxoxHEi8zr
sX/pGednCgB3aLxJp8uU5kSGXfHeib4DpODx/eR+vzWJABYtVTx6ZZ1ULH6lmH74kUTntbu+RlSP
F+Qu6lL0cRNSQP4KtUz6Pw3hU5dlDzITY4lZmUdzzUbR5a0D9LeCdTZoHX4UKyXxdf1rOFO2WSdR
ZLII97GWPDpDK7ryvHPnRYV/K/DNBgkxNPuQd9kNTIwo2aELTI6uu5f7XE3636K5F0qRjWmj5bwx
gQ5KQABZGoqBBAcSMZpJcWiIdenSZ3AwnOZeRCj/4wZMi0LpszpaIHSMPGZD+oOZ4Ok7FjeQZK/m
a45b1FhPw/D8wrccwhYhcdo4CeIROqZ8azNy+5XtQI6xNfhNSPTXsB0q0YIdfPAsKPoRM7FBk8dz
n7JkpWNz3C1gepWHYZSJs9fB1y5owP2kxfyvM0MgZhuEsAyd+WGUvsLdvD3ZkdoWmkgzLVXgfVsM
gMBMbWw8eDM500R+jeJjYjm6fzQOueacx4fPI7RT+rII5tEbYGlOCjMy0gOkKM6ePnPqy/GdZ3bn
L4WXIj4ZjXraZ+Ij5q+ABQVuWcSB1oDlWuZUNJYlAD+heK2N/ZK7+YhvbALd+9SjbBa3XU6mmocH
Ri39ybF0e8LxmFgC8pnXZ1giO+SaxhdUJraN1z2UjhhPBgA1xvg1vH3BGOyxPp7v+UwGZDk+znly
kSQ47gtqo8DKS7GAhCZsmZKE6I0OO3sBwaDENnr3ReGmupkSAXaNBFOXqvuBPwnnnnEe1pMIffGV
6DawSbkOcF1qqGi9vNToz+Lzc2a6eiYDI3ByULvY8iOG2Uuc2If2FT96hYcfVOLG0XP/Tlme8Wo+
+Z96EaRl6PCCRiSIp/xrQdIKZkRXhAMlhJlr/9W9lwMO0Kw5QUcpron3J5dfGJ1SnFJCXuK/5Xlj
I7YuivK7gGRQVQdZz4nF+9sHCA290fA4cYLoB0Ggx57wNm2U35aQ7Am1SWopbGEOYA2y9+9E4ETi
XUetfxQ32FmxvPO89j0gCYTN/809PfdPcDl35OHwYd8fDx2WVRCdpLn5L8j+B6BuxQTbuRBV9ZVT
QUF/BT5ndQfxqnW4NbgmRr0WV5A7Yn/YbR7VjwqAOPLtMo0MRB/U8C9LBgvCzT/PWgfn4YYMobwO
Oa3obLq/WhK3hbNyH5TG+fjaNoEBQapWdA/qrQAOwmrWr03HkIiG+VHOcbh5Rg1lekUffVzCELLM
2koUSQgu/dOfJBNLLqdMfJ8lJK2bOCXHuOZK+6Crs+Tkb8XEp816xHpvknuS7xnRCzye+YvrhzVY
7f6EplkDYXFjX8YqmgbuETqn09gAGNnzceOoA+I/dykmYl6Rd50X0RyvXn/eLLbjkrNXIskbduhf
CkyAnEXOZvL6C0YvSxxOWTpMex07vQLuMUoOfzhPF9sHja8dQeOwNDPcHOAVwWFHSS7OfW/vQwSb
hktXneoIz/McE+Lq03hV5E4tXfujFhf8sPmeVg/c5kPCe8n0aENF1UtiHTPpPjJ3cw+LtGRTvR55
aRvSzH+oINPQgYVQcllu+KQlxysAWxHxdTaPCpGltKADrmh9uCk8nL93/FwunaRubxp+cL770vvR
TL9fGJdvHQhsMPdjfpcBlOGOmMKJQC66/QXVSxoYCpuAe7XLY8c3BSAmOlZecwkGPHp8UeGd7osS
r4kXFexysfQ0nrETUo0y/SDoeTgNgYxQFJnNxmV0O1SHcdAFdo7Pynl+gcJErbJudaOLSb1qWGzq
Na6vlNicyTG4AZETrUpUkfQYUz6TjvZhMlBQbqBXQdXOO5XYH3NdHQrCD5LUGBfQ+2I0eP51ScbE
+2gH+oCVraqiDyvoEjAO2XQmBG/iRfYf+UUoUWe10tp9zTHv2TWSQ9hM7O28u4WLiH+rlcGHCKtr
BO7hR4Hnsk7ZyCCMksuEdqnTmjT28spIev/GBtRt+v8oq7CeLmv9RW3I5QTHSo15iJiG34jZra9/
WH1BJFlZu03gpogTVyRkXHtTtojswZBhXay8R8Ii7vbNvK+1sOhYgXwUc5uKWbWw2MSQ79ivIr/1
hnr10ln+X2Y8VsM8DWFtdkE7j+CD4M1OlCXqCKYUsgTei09kEmlbRuVB9LIXX9wEgf5hUWtxCwKs
212ErVLUg5qtfe3Z/hWZ3gIkzJDu6vZaEBhOHyI0dZ1ZVoJk8J0PbVPg1nXBQgQphcz8WjzTiTrv
UHD6g0RA1nYBihaLBCvRFCnBodG5SN3PbGp7s0LXB9wYTsqbilT5jUorTPXhE0wys3yIE18AyH+D
TOir8k4Ygfmik7zbKfXkbqGWMP3eYpME0kOVdjWRez9RJxSBFkZ3ZryQWCiVIomPW24by5FA7eh6
jjcC9kFoEeNYwLUxObKInTMJUYmKR2z0gLtLmMC11Y0ieor88/YzDXmTL4S2gxBjlqw98mWyeQyH
E2dsdCnNc1MYoN/3gnDW/XwjlfsJ//dQ6iqy/GY+yZlVamH54cS1AGVXs0MWs/9y3UqNMZ+HKnns
vWCeKTtuZJqgaiC1Mmw4QDcVrn2cUWtJcVKVrIY4W0cjN2BEYg8iNIjq/3lV+071mopc3X3RYDXm
enJf5IlGYCyzTBIat+dKkta3GYqXmri/125kwq5PFpcebPXT2nRtPD+37gDfdh1lkL9CORP0zxCq
2/+S5DmP3ZSe5lYlG22XBeGTb97MiKy7VvFXM+uc4XE0t3RMjOsfo8xw2FRYSFZUrLhDEajvcBRW
eSNPzFMn6jTRRhdzFMK8ovIy6t2QN5k8sNxr58WO9ygEiZ+XppfmXTv4g73Ofu9FTchCvrX2T7ZC
IeKw/ghxdmIT1vGjM4Ab2psaatCRTjQQEZ/zOfSBMhQaSIm7ybHF6vl2goErCPy7ldDJKeADbPVV
hhn3rzQT6BVQ6eLXT+58wegEDrCc1OlqwrG+I3MKpJbeUsASyJLYkh1DXl7oq9Op02nWc1SaFElY
XEFZMwGDZwCkfhMAnwGM8DYiNcL4vF7Qinc/sYTGR+gXn3PgIvl9kc6xgnott1som+0qqOFH3dJ1
79Q180phRebTqUGoKBru/5e1qAZZkS+Lzpf8FSJpNLZAnmdHhv4/lwj+VePjMSH2ixWVPnGyaMOH
eueMcWEl6Di79DyHxATfjzbrRbt0LjH7mRgsVspxiS9N9rTdcdih1XgKdN9Dhvc++cxlwizFlTrw
PDtyzk8UGHOU3DoXs3Npk/xWlaFY4EsfF00bs1TuoyX8AoC1gk1dNP+BYA/LinqMx9JN2xVXHzFc
I/ytpJW/ckeBG7dK2qEVCHKCHMCvFqng/KnJkFlhQwphML46+jbvDDW/WxI/UJBYn2vfFybu4AJd
s5f/am7v5iUMdW+ZFHNjfwqRB4Us9HiZVC1AtBPNASQv7FlCPhtiuUec3fvtWpE5rL5/mfkFp0x+
T9tQDbXMp5tKFMid8Ls2jUKofjtglpWfi0Zi4iCjovMHPZnuDuDcZRykbZXKEq5WIZCPKGwM4O5Z
w+oPYRLpX1qnpGj9Q5dbxdgeYPi/LlOpEEjZeMi0AVNumTD/UkDb3VuA7EBzl966IaiVTdMXoxu/
4QmfDyEir70c3kSqRS9ZuAPJGgbDeYrtH6ng0b0FLK63hYCcCPzbgmgqyrpiBkS0K9ZiDNteDoZP
0eehloxsAniLi+UlNBVQTtGR11WjtFQVD58VH/ENxuI3mKisV5jSSgAzMUXRfPpoD1QJeiSwkpvZ
t/U6+EFIe1pL7zLFaoQUyjvO+DNj60ijI9ruAcifsTnQOJWd8D5ywcE/dCw5d6f270iyYFdqBxCG
ZK5EP+HZRtf9rJLPD/3l10KLZCmkSexUDWWs5VaTkclA8p3dJSu/NhA6yFZsolv/oka66XqW8d5Q
KmGXdAXYyCIlAKtkWGRB/JkL3TECbkmy2VhVPOSkVhkgdL+lNQa/fcph/Wd04RUwOBGJqLxNqTyI
AI1ouDHYaifr4i0rzNA/PyO6gWtAPmnSGxyLmW4izutLjkokujujknfHFqZC594ZiDtcO6cEQA15
HPgbPXtwlWae61xTf4r31YKefKD/F5OYnfdTdS8l/C1dIIqNXT2YwEXKpCYbv++AGNKD3Ezgx+Zl
or/sX2vx6M6vplmo2CXb9Udk+bWnVogZkh1eRYTozhig5cj3w+1HwvDoqIo1IpEGd64Vl6XFlZBU
xfpZn/QgOYH/3dGILj7LW7veHfTwZjX2ogb6xDJb0DM9v+k5n6vfOi8iJ2YXf+ORO3SMNVZWNu8I
iTCk8N3nCqxqGXY9/3TY+nsVa6JoKbBGZXpHaBkL5kJUjOI78p2b9lYeJwhaHrFv4XG2W8xo5e23
HER8BYpxB2x4j2j1AaEV3S2MO8ldT85lJyloN+NJwjJUeIDbTw+SjM3UETgLIt5GeEKN3Wq5zL1/
LUEhkqAFadvhRF1QwaNNbhFRuW0sb3OaG3sIXyfXt6aXaAxoAVaWKEfcZwrEfqeKbZfa20RndKGZ
smQfVk4BEPdszQganivpwQHGCC09myVQ/f0qoV3Fb5MXc6Q09FVdg9EUK+XvoEiDlnjqvDpvJOXX
UwBbdJiLrTel6FGTgsMoKtNLKQNPRM8g28R6jQRLcelv1i+i+eCvYYFihAOUlp2M///pEOew6v0A
/LBD2pf4Bed8vdiD7ezZcJwlSCfYfKW5zdbbcvEPrN6OEM1j5hOAsCHvP5Zd3iVJtuB2B4FuWeZb
oL9kfwTP9G/WGQ5N8iM0vPa6CudR1WomIEbTkDoSUTJOoaCuGGEB9yJ7uX2aG8k/ke6RbVDS5eEV
zclKHtecMC/XZblRkQSpVHnucoEVaV6PitynF9lAyZtn0kvS5r6uaPeB1XY9oQA8wpJC2EZPD0lZ
1Fn7jSVkaYg9Rjj2dd88cCXEsmapYabaDzgT/cy7/FNSNow5vuuUISrQOOdSGUJ44Bju2PIdxOVJ
lUtM7o821QDA/W5WpnDodmR7DyiRrGW6aQK/00PA9thW011zS1vFLeNWBlcOw3EIylbtPiVCUfok
GmJCkZyU6/x4h0gWptuaU58xwe6DEJER2dHFN8ZsDXOMGiNt7IdSObhNdgGY5f3+h0PZq3SUY1Ao
/Ey+/vjPRFmkFlM69qktwG85yr6fKWoX8TvtJySmZu3mygWZkta4aiAcXHxBDQoLZctDKb6cs296
FfuG3gOLlwxX/tnttuoeHCV5qZ4Xk4f0taRZShOnIW9xngMYx2cJMyiL9vzuSSFW56LhDB+SIaO5
SLQ15jZ/QGoWnm5rD+b9M+S+tcN5OXAjiqQHk6zlcfgSS743WjLaB1uj9GpvimNKOZIwwoeEQoTs
hcVoDzIWyUSDjY6cyNRvuVkz7FBmS0t7Kzj84MCmL1x6x+PNTi3jGXnxtRuZ0tgzDY9qWK5tHM9o
leKQeqm9yhoMKXpZEw+HYtrg7JPjzo0NDim4QawEZUIPJiHsOSA6Pe/iVZ3+C+1dqpsleq3CVQpi
tnBM+cTKFFXY75wUCbv3kmxmatzbDldsnQXBohlcJPXY8n/AKaC0NXr54a1AgCrXKPUBf0YWaixh
mXm8k8PjuDcGQsDTtxaeXqRoIc9P0SIdVZgbpRr8IxvDp8iJfosW/MLx0IP42FpUgs5vnLEFrYFV
9692oTPWeQvbVAsz2V8WdO/nXd5AcC9d3DILLmCVpiCASKLtgEgRiM32ZVfyGvgK7CYwwmWVrbm3
N3ZXxBuRO2cTY+RsJBrKwbpoWvrf0+6tyOsa29Tpv3OG9iIQpH4qThNmh/jVt5tvL4Q2U6yNgxrJ
Ol1qSLpVqQXBZ23nhzjjaUboQuFBZV6l256Q5w9sKr7sj0GbcygNsm+Cprmllt0AHz/GNBNM8BAu
nrDneLXpWORWZB0ilZk6cxsfGSe+eQYYXOMja1xD2Jx3cOM4h/q4cZLdfKnvYUQpaBRm/r5NO6/2
IDdL2SLbAA6ExSdD2DQ0BGcN0/+2UA+lfk3F9tMGMMS12TgevTFhTM4GB2j/0tQQA3jmfXZGAYmw
d1meOggTmFbXv+l0adU4bzB5EbSqKVSdRgLF87aIEXFElzw14YIgUu+mRT3yVWveaKLMrcbh8Kbh
lUjpME44clZuZRNjDI1SEoK88/KV8+N8UZdIl/7t0jbYPnookZO3rY4NTR7lmV4URnstoSb0BK+b
Mg7bDlLs4f/Du3V3ecaYLzJuxT5C0VJrwJOpgBdN3G774Wxs3JnOec4KCboCHNV3I4btEyhPqQ4p
xOUgE+8/GBtOrwQ9K7CqAID+1jjS+/7/FWv2o0ksDj6sBcXDJSzD2RiEDtJndBrhfZFI1G1t315c
F63sA+WGBSPx8bGUE30qYhq95SDYqhH+HJnL4XML12Tc9QaosxeehOM9LnCJNcFytG5K4QuV00H/
EHVAIUyz6cFt5PR25Djz9f+cXSSgg6sJf55uTCgnJmWk/+4RouICN+erQ/9dy4x/wvZk+dqJQ632
VZKBMupyR6JKhtlwmOv8wtREBoAGi/EQZUaII87clSIAp19EOt/gZ7kYKnDtDVhDW2z5Y4GfP8Wg
eF3guQAARL9AGHKiMVaqzjK7T4nKvcGDRRprcX2Mn+oV1Xmrhdr0Y0rz+Tz/gKTbI+YW9x1i9ijg
IMFlKxUzs9KUixwvb/wQAckcfHcWWFTbjihIVpSVec3J37KUwAA1fp8obMP+k6LjrYDAUDvA6oeg
XKYCcr3HyB2IFc3Yr2Nam0KOBcLDIRe+i6ftr9mHRT/PKdZcsUmodrr5sBVPh1mac1p5YfQA3koF
hBxd4wG6mhzn777Qhcn3ANkC00jcrGVgmhdEcsli2JR/cl+D7E8Xm8BDtSxDrGkPAX2SqSyIxs54
Vne+qCkkhfTqgDIFoZpr/4GBB5qTWL2OOTCcoakbaEUL2Mya8lcBI7lK/yKfj07dEj6alcg6oyE5
RIUdZJp9SV+VuX0rHpYkNnbHB2sNNeTon70fIMGaQYOOULPYgwka76Oi3v/J8VE5ms/dfRpmgHrR
jiMWLQsUBW+kZoE/ONj0hYMFKHgvZC6IcS4tFktu8zVvBWwHRwinQUC52sBrpoAgCgw/dW2ogduj
eYXbwPkbYhXAG6sGSMX5ShSsKd7QY01ZqgwKRCqG/7QQvUDUqndHbiZFoR5l3qnMM5NPqfluKKX7
6EOJaBInPJTHSuWqlc88xId/Pk9AGJKiiOLNlv8ANa6eTJ/6ZkikXyjXT6wY39pfd6yIpy5JYc8+
S8zzLJTf6BDMv/h9oJ61vlF8qthI7YnKNc0LtcYgC656VxHekzh4Y5MgHBLF6VS/IWQOBgOX97NM
Lb4zBW+HBFVERzx2JZFoy3ul8kAubQiEZA1DR+U89U9qbFcz7WXrcT380LMyY5vi5qN6ysPYzeJV
MFzGLE33gjG+7J38L/r7IERgPulTH3V3nv6vYELk2gks1HIW7NXCYz8FFdpB8qONRI+esnKIttGI
snipvcjhhDwm8y0g9DleLsYp68DKpeut6yPfikTUYAIAlHbukDPycvhJm7eZXujHcvvkrqkfGOjf
rb8HKKGfo0SxkpnACkoBLEyEdF+y5G4/aPtEOZDjssVv1jjhn5vD6VzZyZBe4fhHfHXdqBOA8mU3
gOxg0prPXczDDYOY9OSw8xcrP4UGidO7gDRIVnmNIspTF4W+/DwvVvgceR8u7XMcQUhQcMctVeY2
W4bWCqAq2yDTHiZ9ugPCp8b8AqU7Q4aJ7uwiYVYaDzH4fZwQSt18miB9AhbEh0BEvBeghyb1Rl87
7R9pwT+kkz5oeEd99Tc3rxpUl9ZQC5XI8Ki7ItChU63DdsHN3v3luRn8P+af1TVBPZNDy2nQXuwd
5V2qLpoiY31oG6QA5voONUihguLRNYavFFXmlSauDlaD4MyatV6FH0N6Ir9+T/qGt+Qn/R2/8X/t
ICmn5g44E86X/LMD4j4MTBxFh3qei92kLI5lxQWcZGqbu0axWaG2dtoavNJit34pVjOOBsPuR3Vh
tTmpC6XoTH2gbYDy/SmIvLidtiIj7S5MQzpX/t7BsDfSpYn8ROiqtjjYXdKcqO/OyiCkkjCAX/Zh
v2FnfXYu6ilT2l/wcDmB3E3UbuSpsLarVkX5zsnY/gF9EXW8G145PIn246f6426KVTh8EYSdXdLV
Mvw1DQR7w0whvnPA4llfKVjPmiP8rhilCplwJGi1muQD+8bWBtc72F1NAiUeTRG/JVN/pJqryXbr
bz5veu+xqtYiczsN9+Yd5GDr8EORJEOeCgmwovQQJASw96ySKk+OT+v+4zLgo2qpzx9X7DV6fY5y
6jQCheYaoxmgK9RhNsUPdwfxn5j3Cxsaly15iJ0rtyBnbYnij7Px0Edi8Lxseyed6/i/ngmn+9GY
CEnOQbfYnVjLPhOJKOagqUzc4/FM3XzgOgZ7m96ly2W+KU2fh4znK78TokiInsigEY3rdq7uaRsg
mwmhvnlApe8EKoyM0dPDh8THU/9CyNHJoaLLOk42bg/VB8jWu/cGzlrmatZD8tccn2FcIKQCdMlT
r9+ZvAMtss3a4KQKOOjnIT7kdCKk7ghmS5S/GQSlb3LkeeRZiKAWkMKZSMv9IlWhUtJzI3N/CN17
4jBVS9rEZIujkg/VNnHDmvQnX8o1eQwrlIhEZafApA0asskAoVZ0f0qSfskTNGjEsZP9lbwlms3j
Xg6GhAEqhi1/+hIB0cWaeBVy2axM3z8HVKYkUIy1TEMRHOgzJspcn8GH6IFO89vk7q0ZkTBQWAGP
y8w7lo8vV1Q789AFpv5uwDh2HwaZBqJ84m5X/NqDgAf23ZrPyOPTUMAS/zGBwGn16+7ySf7Qp6Yt
f4AMbQy8zS4qr7tY9fCRQdd5gReHITfu2KDSrAzGMk0Q0YI4fZsPkNQlbq37f1f5KDdrJruKmqvS
b2Ma5g1K0g6fxWMOFcZ7mN7psyndv/Sdxj1xg31OI/JVWv9kd7Kj5ObSdGoP/9hxQPDJAFq/Asqs
jmoiuk1p8gZep99zX2SfTjOyn2tr/Cghkd5EpyoozyaKeWQZTi3Rhb5nUv7FsHJP4mqlmq9ZxpUF
ARRqpKWZ5/Ht8ve9o4UrD+RIl8pOaCgwDOenijTCqrZo9mdTnB/Eodqd0hNJ0lqh2J4CRqyHeCVi
qH1xptaa2tnZbmluzgASHtSqqQOf1p1HBmWGTdNc9YlQmtnnsUivcddzFzimpCOZfQue8rYX28Z+
38z+7snH5o0ecPxYwk6MKq5377dPJDbK1VuFudnSRaxMzKdrGOdVPaowGxXIncLgdbkoNmQUmm1P
bAfgFvmp71EaWXUYGvrTT1vGwybzPWX0eAfz/xjRCF2OnybElHY3HcXNVLKoEidvcW/WXDUByaoa
PwhHvscGQK+4XY+vt0/aORMSSkXK/PovqQYtboTS0QJwDtN+orPjqym28JM8wEvKrpvZE8ZhMHW+
LvholNWSp2thshyZlTMRBemPCfKORSd4eprS+gm+EJM3Bxs1AjvqbqL0LC5adlCeF4uwFDWaYlIn
1Yj7TVQQJNpAFzjk2scswYjyIMhG/lqR7Yn2F9QQP3Joq/1RqEi1sd+hRkVyxAJJivtctuGqT7u2
89XSkfm23IP2SiYRVydke2q+MfFDnvXvBdFARFgCCWZbAh/SixPsLs4QStnj8DyB/xpIbMzZzNSR
D3/1q+7y5dLwu07EMhpG/hnCj/a7GLuGpSqLJP8voGV/HMmYwlTt6I90SB6QrxCiH/ziAFOFLW84
fTWLUzDWjI4OkSwcVy/86vebn4gSGMxx7ZYsmZ89PPQScMpwURLkLKFTWCFt/9dKVeotM4LuQCaP
As2dSev2jMYDN+kS7viKWCN7D31SQ0OzKnSotW5FnWcU6tDkDLGveq4fTaKGVStZiXBWk3O9JmYY
+Lm0+5Ufv51DPMUuo54LQwwzYRg3c0TCscbpiIMxLiU7zDUtojFjb2PMGvplHFvR+GB6c2WkLd/u
5cgsNPadq7G7OswdFpsRwnJ6wY/QvJYDE7WyjoPMD0Qvz/H4N1ITmCsz7wU3JHIG3WqARR4cCiWl
3xDlJJ7AuyBy3MdLagykGPNakSWZAjiSzwYLF2pK2Vq005fsYl7Iwp7T7g43wSUcmH2HgRXpZpVg
MIHZhatR7bt09aPnA2yhefe66ZZhb8X4cvfhkwIG1baREejvDYtriincZQhkON8F43tUE8EJWfUO
i4kelNTYqFUo/9EgXUf8I2MZG5Wroi8RKnYKEwYKn3kh+CRP6y6YryIF/SkCmRNacZd0KmOesFf3
/mmeJFbKY59eyAnE4pZjEModwItSASqLpTmhD5RKUvJOBjHGGlK6xVi3+I8P7FqaUQh0RQDB43Fs
uWbHajTOXRY476ZGKi0kmvwqUoUVhtxpnJHYaqbveejsT7zGp1SULGraE3H3MJNtq8qG6ap8pMvm
7JejBFz0AfMq+tiRaXDuf4F/S32hGYGAAIwT5O5ItyARsJGWbdfy0wYbUE3zfU0Jz6htf34klq9v
K6jKX9FRkBmrRJvfM3QJCyyXlHn2gAfABGL9OzBa0nJHa+yVjWE+tO0ArXa9BFpZW+SUpmhET36e
u4rUM++9PtubhtageRDlpnn6yliOaeibYKIpduH8hn0pIcRracr4dCVjjpm3pzCiLS4cwNNLYZzw
KSP+TZ1sBb3oUZQLsPplR/cy25jopaWJBpzdbslT1l73QMw6ITvqH5JDhkzHfK53+gG7X0kfHdaf
hl2uBqzj1V4cujR02bbJ6uy68vetrkt1ZIBQ7wfj3IxltIz3geiOaTpxlmx0l7KeIvJkonsr1qZj
jAAj2ijA65RSXzJ044megDMiiPdyD55gubZSBZ+RGFnLMosVDsSa+fDSLm1QfyKIkO3Cs0maECAn
1+wGmxKX5QK2IXkMcmpvK/wZ4Dmedt2qTGL/opJPSLWOwUcWMFWcgotykFnnXPsnk5tm8yiX/dRn
Vk3+zfuYYQZ8ewTcLTxXDUZ9tgVuZiZglu5MzojWRgD2WRAhY7FQYefCrjXHcXBEwO4wwOP0ytaL
YM++2BF2q52Wv6R970c5GXEiuBxjSH0+NhfC+3RTc6/VtECKX+LSslV7wk6WtKi1gVdO10u9LAEj
PG5gX5+eWvQ8zrgdXNqx4/e0bcJnHzy56CZd28iOLuSnFUe7kiy4M+VSRps7Bwy9kYl75m+T+RFw
iP0ez9dc5aX3ft14zSSIU13O4HBDAJa1h+8py6PQpyo+NHbbTjI4goIju6LIxQBKtgDJYrqHTc+Y
1NsLcYQYrTXCF2guY8Z+ku41ugHYDog4/vHG2EkuSQqcgojxPsiudatLjJXbnK+8pyBkf5MOsO22
rowoe3pyiaMljhDWNc3Bnk3ScvMpIRCi1G/4AdaXo+AeTkivI8IE4CoEmINLvAI8K6l2uKF0XNJ1
W4/gZ+yrJqv6wQ+VG7/9D1dGrcd+RDiyGc8vDNycNKnynuPUlYPsrexu2svm0QNt4TIkvzK+5TI1
NZmOYATcsd3UQokJHJnYXTxVGSkxa63hrM4IP+v1tpFfVQqnzJ1Rs3czhKUngNMmY5B7he8QTY55
40icom0X0WsBo6HIYmdBhkUY+wQQrF3bBpFKCKhnlxekSQwkFljlIjNqD45XEbhcxJZXfAw+pYjv
kCSJ8/hALNOnrdpb/64xLSXvYS7yRFtTNArEvNSU0nV+2ouFkU/hB0w+nR63hp3b+HoId/AGGYpc
7W4LkMoLrb63Kv19/0wnlsGJIS8KODnf6WYIC8R0fksxAQHeOk2aude86EbEttlfNz/oh8DcF4/c
oZZdKOMYEPfY5k6mgDwA3fsZ2F76MrDYH+cBvjece+F5VJsoYu7Pb2NRvB1k5iXuYR+G+1iaoCcH
+M0wSKSntb4qzrO8fjWZak96qNlY9w60BBmOiI/In9TXRtUsNlcxRLLLmBdcYGCRP1CyxhnSLvLk
o6Lob3QgUdHkwH4Pa/++5y7jexYSKpy1AznmbGyGRxf6H+k+6dKABtZivcpAstVAk9EF7s1BUeL/
whxdqvbje41d4j4BaOoxrtWcxcgQrgpJaZqXvfF6GfZtekft6uG8CbHC9acjqcYh/gVOOHS+QF/6
C9DC8q4quEzDYs1WHSLMGu6o53mrI0MD72aQPd5G8Nb20GbO0XrzxlizWa4TYtASgHW79ACTGl0a
oPfG47QSkVCNBjgmfyUq7iN8bx1KMo++So/sFCmy5hARlZZg8aELO6SnhsGPlxLrcWySSex5NJTF
wrMOXrYRwxLURfteS0kKVgmLEn/lpxPxyWoKXppLMDfIZJTs5D2yHHB+ApYROeIK26p/OihZB9a9
hvDz1zVXFXIqZVmXUIpV6emjMfre3qfnjq2CfO/Mmri8isIHS6IHDTh5mXGHb9E8jRQPyDutKoLw
uOS85LDtuqsZeOXhvdeUncmVYLwwc8nz4SFrUwgZV3KNBMzi48tJEtBJSgcdua7aSjzQqY5CJXlt
yqyi3Acggg3bCdbsf1upzMnKtGhFxC+tqj+zksaw07adGzkKgJUowy8+q67tib9vRrk20PoNIxYV
lcmqLAtvWsqOfchaTcJEMT6ckioeY0HUwlc383gI5Wqm6qh0h3q8IRWZlHwutTnVRkMyxFQmYRS9
5rndM7uaZ1oGAQYgmwO4zZqRg2WM2PzcySW4WJQ3r/DUB2UnXDDHLkAGJqQvUT+Ka/yH/3ZvdXLm
4U26LENrWnd/Hq1Iv57w8q5+NxRXYqAAJ8TFlcVmdI1WK0qrGigKlvMdLaS5jADpxkATjqVv+sA9
hf/j43qTxsjTnkeqSRQT77hX/sMBcD155nWe7wll10SWgZis622d280nLsoioPS1IpoxhOCd+TpH
Drur52AjpqX8fUEXxhVwxf3NrWa4SVqEikH1guOG0AGt7D+L40h3JxGjtVU9c2RBawBWIwPVZ2R7
KMmhrACvjAMs8dN0uKIR2OdxB19/pJIL4qLqxbwFwUza/Tb8MeejjOHQ/6UaJHm0VekwoAaYw3Pd
KaM2rA1GJzFxAskqWwjO7em+cODfiR13IHswfJrt59tMq+MP8pkqnFpsx8U9lMmHPL47+OJ3vdE0
jF7pPJ0OUMDTbAo/2ByyfDfuGLKB7VbROCaJDUSdLPPgtQc236bQYUmV8M232iNR0BGDVkJdcqiz
mmccSFZG6zJWaskUag1zn57tBSdKXxvDmmvaaip0lYNMsSXLLQdu/vQiz0Qs5TYV5adxtty++wLi
5v7OiHkCSrpZWbQI9bX5d8r6BKq+DAq6Izq/qPZNegIWFbL2NuwWCwl5Itd0HJ5UdeBhqBAxaz1M
ujtR6o0d6qYyY/RiBNXfbFywIn5P+Cnv+aCRQCB0ayaCCt7jyqRHaUBqrFsHfQNTqW0f7vZrwUO/
v3kvp7TUakmEw2D9Iw9iQEU4CCJ8jTpUUFN2GTpx2tWSjfdLDdkizYtUGrjZ2eoRVhPs1lv8W+F3
AiOPdqAW4sEUeaIbqpq8wN4YhBw9/B2VOa6rGMFocPZbxqEv9qbH6NFQ1v77dXmcO4qa7nqSnivZ
Es7qQFtgujUAYofnHiVmZ0yQbrKsy821Hd6s8NUaWF+8yYYBLTIr0wA4DQ626E4/zme86MA8TkL5
YJ2Mgu3+Dw2Ny/eqLIjXlrOMUJzsOA8VA+wfI1bWW8jl9T8bNDOKg9+9rWGGJrzPVF04zipCSQJ7
IVFMxydGPMoBDEBaCMP9MgTGcz6oztkEVqzPid/1xeahoec1NthQ/tI5Q6dGlsGHQlcC+VV6Hbx4
2H/YIARimbq84iiaWFVtfO3D3HJ0mIYrTt42HAypRW8NmFQEZRyANcdB5U52hjIrySnJZ1S9npp3
ghvIVK5714L8xKra6KCv7ZubEmx93K/F7AF+99Y017yczhjrcdv8mTbKVWyvPQfG9cifIUcGoUrx
jJ1HTkd2vda18amOSrZH3OxcVj9REUvHYV06qIJeEKAddA538XGEz3ICUuYB8pxvNEufzUZuIPC3
WqvCV/yfzNWN09NP3TydPxdB9jwA+hN9tnaYP4xyBIcW0B2CnA/1LYIBi6AOKQ34lIpkccrOTYSd
4CnwlZ4MBxriI2tSFj6muilqeoRRcayAjOXcFwN0aq5xrvyKJb8J1li4j2OBLdrY7eAntvjB80ps
EWpxPydrW4xs9L0MNkAKrUzM3IXnyZE0gKbJRCcwsYNidQOtJ6ejYlGvzUY6Sp4pfEvDZj2P0YZN
RHpm5zeDR/qxvICofg7QFuKVa+ksR6hFEa8v3eDNaY8MXtfb00AU7fGuKcJuWptpFMVUhVC2mhFX
YcJFstV9eyPwiWKU5f+gMIE9IMZXlkDtCTBR0yoJ/+fsYZs/8qImtqeKNLrMyQ8xroogOzUjBXqT
J02UBiH5Fjnb1XD1tGJF2E0Dgb7BCjkIWtvqKpoy2z1xh9Hn7AFJSPp+8UV0rLDvItqg3WWOPKr+
P3hVPhpG8Ehi1gcYs66pPEmRRanR0NUReri9q1xMFDALBbTZySdIecTg/HebuPCYFNYYetpunKuz
ARRPoDiXuYzCieMwyWxlhOIbxGrJAUmArn7B3vUQ5BoUfA/un6mi9qBSfgTZU9aOkmtwwqypnCtB
A0KdfJquNJCCycMbLZTiNT9GQGYqzQqqAy2+PXdVQYciZrCnZ7nLqb4PMGTdV9wemxmZOEQ/ynwJ
g7r1OL5+f/S/azjZlkzM4p2FdUre/vV10+E0JiRnB7DCobqkrUUcZfsTZQ8dN/KARKeUP/WiXcJ+
Z4Onpk4edKIj9nqBhH0Rvrxu49RNs/OeV/8HsqrbvT8svr6h9QtfkaUQ6ktrXVdzZCkNrMfANREN
F+07j8o2iBjaWtL0pUbrC18BwQS/sKfwvARGSndD3GOnyh1iUkdJbTIEx8Zs90fP2GPqq5FxGlQp
JtseHEAaXHeZ/sW5BJp+kXw0Rl+4aQyuT+yiPg9Ic/1oIKUD0GBYtPiTzClgon9DnH5wd1KFSZ+y
UAoKoiW+1en/K9Ysp+I8ZXeZUNnMUwLwGRbn0EFDWSHVxCRzAE315TY3bz9+X4W4I4AwSTPL8xZK
je2R/HeTkTmc47+cDDvbqigXMyloXiM6xQ1gBjydDU3bGh+tuPoyG+d+Jz7J3ggeolSkvpS58Z8y
TeQ5g134SSz+FsEtBcB2bPWpg+Gm4OedHtaTn97vY9VYmAU5xJ03Xi38YeuRUeMxwzuZtZQghMB+
I7RY2Q4qr11IUDFvSuy8I8chMa95LT/fgs4jj1n1JNTjiGIgNRmkiL3QqTf67fOY2o+0HMtO8nrU
36zrCNwjY/J+zeN4X/vXAG6uvyBbMC1L1Rnlwq7TR6VeWM8+bZo7JIcXmbKHqsms1pq5RMYTTaAD
j8mrDP2h3iUEA7LO2Y3I6YKYUYqJnnb5+13Dtiacba04fx0dhVMxlMtPsIPNqAj8mczFUtaSi5FW
OG/Ds4eapuk+wPQlOfGDI/I++yjLT5ywD0R3p8zryOTpJBRzGt1X71EkHqxY1SG9Nm6Mu0rkVDaU
Q8Iur608YOpluSrIjlqzNJ4r6DiFTN1YYzrA7ePO8F8Bi2gqDdPt9ygqtrKs7kWAcF4/x+34Ri/f
iaGfd6b3IejqE7JR5M5ppzfmao/7PugiqjhYXPLy87CrqJ/daQIss3hSdSQZ0KDX/7Sh5Pt3yg1W
aVjxbFk5OugRL6BP2NonN/F2cXMSu1QvSurP3a58BYmsmqc604jVMuBHyGqeN9MnovZxb10KtsaD
8xQSxkfNxQ3MS2lBD0p7DEcwE7hkRyIhd5XgClfe7xL/m8D8hRiP7k6jvwbVA1AgX8cH16BXPTot
LYBEuuiMobP6mYekPzrReS/Ng8frL4U/gejaFL6ikTSP9Ky8VJDe1RzLQZX/WnasqMA4Aq1TrVoI
g9ikrvCzavS40msC5JxqNpl2eIstOQv/DrBoRzL7qwH/uX7YYvx/J3vwAk2PueZT+zJfHOc+deqJ
Uh9qiUmExgKIPszqFb+UdrvYbJA8Zz7OaU6J408ZrJ/UPI6jTSGXwgchk4kVbW7d/Br1G5HKNS9x
UIilxIX4unC4ZGqJNBGtWvFGSHXU2JjV+KXf9mJHTxJCs28voZ5DjOTtw0PPY5v3oX+Myi6VyDP2
4uVVN5npvAECkf7Pxhh1KSx5UgwZmfhqefKfSM3aa6pPH2Q+RPEiNrPjE+zqbdaTXA04XR1rFL06
TGjrokaejuqDX87zqyon6kLDsAW/WkzBmn9iI6XIDtwUyLY93O+dA4K4kj2ItnLRfSGVaGRBoMh6
r8Do1UPzs1hAAH4kn2nnniCwLwGPTNT3RHXGMAIVLi3PTrUTWB4HV+PGhAVGVqu4ihO5m+VO9tYE
pUgK9nZVTWGr7QuI0R8J5B0FQohoWLOf0JGDq6dOi6B/3vNVSWvGp/jqHZo3Pm9l99iOThC+7TxI
yGk1XkbO7ezib4gX/zCDvb7HUSlberom73fiF7C28avXDYl5/jhav1UZ4hGuZ0Put47NXMbOm3Bi
EOE6cJAZlMezr50Jhvg5eOeeUP6Q7wk6Xo6ar093oQP542O19zIS1lt5a+G8BWmnOJ1zlqvH18Bj
h45giG9m/eXWaNoRbDdAsbo9q8olrl120A45qWlQ6TpkDaA2YLbXXFduXzQu7gdcuETGyjLXeQHf
90QMBNwrqDi9uBSUB5MAZxJQTNi5Slw7UzzH05ek8THvyY3Jclsm72oiQXY0uoD0jRKqBam0+63P
eTxodWYZr6hqs8atlkdzDbcloQGj6HEiVhYA9FCA6ENPYDD9IKjRiCssba4JNkeZWdL/I9HTbzVe
WCNTQl7dFlu1XU/twbwJVsidKCB1mUF2o/99PkXPqb1o18yDHyBialrM67rljzlS2Tflo/ooOZIU
Ng7OfiqcLAu7flND1Nx1PuKp4cYibZ7izn9GRC2o+hB2F81XLwalj0qCdXJ6zYXEWcTO1dK5rzTL
CMmSjfLtzHemjAItGXdKnWqR0zbsriKyVTFe/jJYkvEomUd6qluZhxvxUo4GN/MuwN+REVqrO8Wz
TY5NtdvaMnJnS3ckdbDx1GwAjF9UKN5zGq67jW9J/N13uJFJHwhX5aUQj8qZ603brYq4ukEbJycE
JVoCYReHbbSZD0ylTf8+moxka0u7IWIp6TuZZecR0Ij9+WZv2jReye1+CoOBGCfmJT3B7bg1OycU
7cSDPDQqrPeMUSHdFwsGNPpjWRGHPshonAx5QWSDOjUx9u2z61i9mEdTBLurDBeO3Up7MrOSzoEW
468E6S/5uwrt1sGeO/oRFY1vAtQmSa8/06qtJJaFwd4F49nXjs32mmkDJrYrm513PJCJJS1ppGYj
/0ORwbZt/C7b+dD/hk41Z7d+Cr7uO6kAHSYePI1iUivgDaqI/ycvmiNJsTJP01XtboKzPKfKoSu9
mLYrtU40IDRNc6GtnmgHICvtk1AlC6hSNJKW1QPHaEhUpddoWCoW4+TgneUORsHNAYKL/K+1jVq1
rf3oCfA3HHK3JvfsZtGKaB5y9aWLiy+mJdtJLpHIrV2M/9Jba4fRcacYcakgtNp2T+vOVhioYNx2
77kEQUDdFSUlifwEMHtP9Go0WTPD5s866hupgNjIsAshvIzbFkEvp1/K4gsYF3SXd+7vNRiv9OFG
xXU2OSMeiChF1TFvCY8uKlmQbF19BoaxeK7FTlPJoVNKH4hAH5DtphXmCkB0CCTX7KQaBbr/Mvcj
Zao8+8KrzFf9kSfolm2YxSSlmxXwJLh46/xsCgbgySU4qSoJxvL1mgmy9vsUhMzP6aadeZDise2W
LtOFWBSSXepwBFeZKu47H06CqZ4wxRJzpQ9AWJxaHb3j/8GgdNSZxFEDo+eoUwG12QKn3/DKCCRr
Wnpl/NGO58nx9tWD7pFu19c4gnrKLnR2iB95pYeURYYYqXITYWQnECjIT6204mb5hH72S5uVqihg
2Yji185q4kDFDZU4fdaZ5cjUL0J+biDcHvtZ8bEz8wscmuKYxVBjTVr9dlEghM/W2m5gf8X7S8jA
U9t8R7r4jM567N5CvFC3IzdRw6VOohN/jz1Qf2FnVUhEJDab63tIUi9CpEKpHqrDN93bdsQc2nMc
SHIVzCtTxw2XMVG+uwondeqxDvBjdjwi4rWkP8fDvt4liTqdN6+OnjkhM3FhDfPdFKWXtdt1snJU
vpi2ZC6v+vs2D+zEDncsvJvc7bDBt4qGoySAlj+p56tJ701kM2iX+xlNrZzSJxF3tvxcMKIH5jG8
PSdFRIpZtwka24yGiY84mikbN9z760u1LeRM39GKEUzncV+NNun2tLx+DM+BxNuHmuAoij1a8Luz
yeEUaf0FOqB8veVRCDusuzmWNrSTzTG0seBwzsLxDrl0DCB3YIb7rvivmoaNH2ShbHtgivnJLCJr
hnlLx1WcUC+FgMmRCTlyRWFbaAed+IBAcOyevN40VCt5jJmlYwH9vcfEtQ+EZCtaQ6uDd0E4JVrB
3wUWpHBPS9GzKGbjl0UDp0/fRS5D1VM4qyS3vltfmVntZP1XKhtJMmmCgIYHZKxNAxscInKZoUHG
uX1psJRTAzgpSWDXf/x4HLmpHKa9wZKUPrx86W9Rv72HE1q2FsZEOlSNh8MTJy3rl1DKMgs+Wudt
duQTCo+cCNjo66njJGAS7YGmfqucwdwYJCRbusmzCQM9TXz1+2K3x/yCdGGRTeIXsCjW8hDe3FsW
wa/l1y6aFml0P/o/7QZg1/inA72n78fkHqPhNIssykhuSG7CLivmug17wsy/rcvPmalAuxyItbOr
O18tr8AbOHzi/wSyqGeA9TSyLZ5XApKsmC+zeUONBgz4eeyGaOHj4jOb4MmozzMW6tAV6TmHyNcW
/Cw6g40VyvRNUbVaz5T224XvkdgsA7gKVefxHtE/wSTxdu7CDcx4H6sDzbPCo1faYwOV4AdMJft7
dS93m0vPKMVvhurUR2F5moi+wf/0V2nMEFKffmp9R/xsZ8hFHwE8r74qHVZkz7CuwKvcWFOFBkCs
M8Mem21ZeO1ysBRTuBZR9TBOp3jZ7eOsmBE1TGGMC1IubZQrCNW7BhUUDQIRWi5AhiQIB9uBnzEn
knQLZCwd+ObTHgBZQp2B0RqkFz8vLzvlZMnvdQSGftwXO+BHN1eGwzZCKlbEkHHkJUTkMrLhKYoO
hHLtp8ZiXnG4jzHDcZIpQKAvZygt15wNEd0XmDP/XOHvQ0QDbVg5pSnuMZh8hK1faIFFfrC9pPvq
XQtpa39L0l//EC7BNDde1MxWjXLd5NcJ5F0Eh2SGf35syw/+ZKi4/3WMPFsggIYOGoyJvpgcqqNl
UlkLcCZuuhQMAV0LkgSgoelMUHBTFgPMn06kyBB954q4aa/JGff4oNYlu8d/zdtFeJG5HI3JQJdv
OpPe4LlwhXtRX/pPUcAujTpCTD+bDJFdVhhdtSBN6qGnGs0GrvMYjP/ACu65nMETrIQrgpGIFEl/
CEC2AoHvpuM31A8sBYib7h23PiaYZu7TKzn8J0NcJGAO6StpLNRinzbYfDgFAnS4oPAiCuuMkG3y
gfsrKUHjbou1oAhPUwAmcmIFbSmhm1YSojKkHZxWLLmTdOaEC2xRlXoW9FovlqKxdfWA4HIwXipC
7QdPldv6UgNm47hvTmBDMSKpXnCx0rnHj6VCyRXjwoqT0/m+kYCFrW13hkOAjuOGDzsypNMlB2po
mJBAVLC4ff2orZtHzXdF6XQT9BEVDuT+3n17NkfOdP8TuPKtDIqEbvVmSLc0dgS2pGl7NX3giCX2
iSw945almFXzfw3Vobt6V0m4sCsRV3oRwK+/Ofkd4Nk3WN3emLOCeUzHPXJcBuewz7aGP/+4tgDI
iMVfZiKK5qiBYvFUKqmFZ4PuXjUBvUrNnOtv7Sv22z277XrxhaYewQkSizRGH6AYUG9wuWF3rZjH
spEg7qG7xfl0iyTOKYL5t/CGT4dpbZSImI0WiGatImqBDp48KZ0B5sdtB3nRJmRhwwCue9nTSrau
8hqSABw7bzRNnHg8hFf+Gsm3KuXYhAwOiM4Z/ctuUWipXXnJah3AnrBYgf2skhsWvMEXhShDbBKv
Erb7OQDrlvh1MgxDhPLMQDk7mW4gWqB3H59xuB2ELp3ESUCrxJkTSFhnpKBltkDQ/kg55znl70CB
nWsixmGrKWpwL8xR9AAcmr8SBibr71w82k+4SbrupFsiAdYD3Mo2jzpuYWYlDypiIv8mH2amN3pt
2pJdFZsTYKDsVwriBk0AfFiJvBTf0LpxCVe8m4b/mWzMF0qtb8FEr5yP58ZyrL7nd4Omi5eqRSuY
dtS6wbtkFnVnOfIb4+qGU9/mH7fmxwCQZQW5A7r6yVi21BMjIp+s0eWNxh+JP5cGH7xXJtoWL+VS
mB1PEf2aWBffJm+dVWPNRaBT/FJpcFdZuWq1brWr0BgaiQMkSVI1NCrbTkGFLDiKWc6aYjiMrWdc
AYSaTXseI/U8yj5t6p3MDwk3mkLCEdBaysADmKqHnvlwLRVx22aHpd47MCk5iK0drEFcrpV8xGDp
mQkRfT3aX1QtUjJKsGamL6qR9ejeemYaPkuqrzNeeuaxhIcdKdzFMJfviIlqzwTurSd4idvTwzZX
HvAK6A0Zbq9Y5EDGsJkViiw/uQSybifTNDytQGS8lijTXr2dnyTUQlrxqJpW8FL6P88pkOFz+2B1
v+19IYKorOz/A7RUqLAZ2V6UzHa/j9a2M572YJTN4K9wcNRsaS8ocnUaTj1yhkyBNFoY6sTRCXoL
HHcHipB9DSD8lXXFDP9KjWTXAP6k5pMMXJkWU33QEkB6LAD74S/g5qh+s1qJywGXvPdnR4E9+qRc
VzPhxNp9gGl+V+mfNzLaYkr0muK/ysm/AoqLqLKgXq2YwMsIa7cAWYvBKm1Pje33kxRNNRDbl8Ci
bnytKoutwmBRSRfQG7vm6lloxEeudFnNVPuzWhYTR3n2YB9AKxw0nbO5q4xQWZ/+h3RwLxWxtdj9
cVQ1U6/CQXQD53JJXV+YXRNHmMq3Rg/ur3kpMWjco7TGhl+MJ6jVsVKJnld0glZyOz7Z+/QhcTfy
tgScCTmnD3ChHc0aU+VFBQQhab1j55XgKTSo7e2LnONbMYbOfzPfBtf5dOBzRLYI5PytZ2GL3BiQ
bSHtILWQDGuvNE03m7TJnnO0WEu60Ni9m9mi7q8QmKAv6mMrTUHL/ozw54yab7TE3zHjJc7VIlNY
w6TP3XEgcA8W7f1cAOCAGRGqm6pyYRxkwps2gLP8qK1UfulVIQutAmNvBzRIdLJEWdGyL01N+7ku
Q4B7l5+2qb/6OLcLqtCO1ItxflEhlw1qHm5nwBOq4RHx6cfjVI7ElBU7nP3uTek0fkk+Z8SQCSyA
vusgtQPPuMi8PuNVZvSnDTgX4EZED7wDKM++WSFAetKD+IVQ79gP/eo/xvI1jR3OhYZ+gw2Dl7Cw
MR2Wc31Pig/SXLN6FerEQRTbxJPeV8xTi8m6EpEoy181+9XXxRXrQG4wsX2nkxi5Mh9jdidiyvDm
arQoBEX3xYtxB5w80t+9iFvAS328fUMGydqG+w+XEFmZKjhrAcgAXCaOOfMe4gYl/bh8f3NdTTM5
7iqJXzH/saLxmAe9R17kBANjXGxfxjnSok6vXnegdM9mBAQ8UnsPc3TnDp6P4FpmOX5an1MmW7en
mlNVeMyrwSGnRXuP49mjkpFD5Ssi0i1kq/NGrnyJF8+TE/VmfYomcx3bhaTKwsfUhrEY8GQwdX1K
TfQEXuWtM65Bz3Qm7zV7BPdfTmxBzHB8f2pI3iZtb5y1qCzA5j4MBhP4krKhNsWYEENq+/xJa4H/
GZ//Ev73SDDKEgdY64aMY7hcpU3VxQXx1/agVtE443aGwdMsNRPMUGTu2pCcWk1jo8km7JnKWtvZ
/yA5CGFxKiwqNTnU00JmixkJBYVHHYJ0NnuqsSQPEWZqPiceaiH5W2+U9w7mSKX8JXDRijkXXG3k
1Kwt79BqfdmJ4ksAhVMf3dk1cHNUDlrD6FC6z+AKTAxztairhglCGju/+a5BOJmlFiHi3o2K0ZNj
O+qFpG9VbDq/oxnaxdSnEHzayWBzOT+6zr1HHIDo5miE+wngSkU/KAJIIeSh+r6PJwygrTvCe+3c
XLDfgJWleFnDmLzIl60lXH0SiI5RAGs0IamZX0zIBEbGCbOvz9aFq57453xs1UtMNFWeNw8lmENv
iQ0OsvxMQoeBEVTbZsLBdlpS67IawWGWXQMasOBy5rjayFosnzQxgX2CmIiydLp+8LG2APrI/Noi
wEl1PXGm4k72zQu/jKzgnBPfa6X75+elC7deK/qh40CqjmfGexULNoQLlKD67SqEtcEbYJxHArQA
e8pQs9pAz1beKPlvhX5wIXnEEFVdxnWMA47JTL2Www7pk+Ex23hG0u7DVqBz2whyAhYkhFkSY4XQ
ILUs4d7sUAyNykC3itV4HnNVZhhj5IYZYl2w3/SEpY7EMdxDo4ky7CI22y+PAxFropSgto8h3ZMt
6y8IjGOYc/TRnClrBjrIcR/7s/P+OmotHZjEVu2rnz30NLaKZOmkxHzBZHpF6nhDWBs/m1ixbpx6
tVpNtKSSuK3C82F69mFfnURuIih1RLeLSZVPHPJEGZw7FejFwex0F7kZxmsCh6JWPZJ41wu0eFKz
gpvTfs3VmJ+/szp7pU5kTPNuoXQZ4XmTrqHIvkbx2z1gbwWqQ5fixoEP0aM8iiuyHB17hBz3NoU8
OlPGfvm8QT2QcpFiwAoodQg3j1CVASzWXdEqyT+J/A6Og4xBE8ZcmhdXc3jeTNY9XID0ny+cPSuH
bnbfA8Md5XptE3qPbtYHjqo9pHfpI07ACHb/x99UZ0Z2oJgkCASa0KssuCXJNFKboj3iaUa1wiJq
RlQL9rkmxBDY7o+NAeyKRHVuJNf/7dELr08tFF7mJcKuM9k4CoUUWeGQfl2Q/FDYhNetr24V7LxG
yni6Pq7c7mvw+jb3sJMwCJODPtw4j5qUDTWeHXfb+XEKedj8/nm5xWZEWTDVoe+pj97XmqIwOBqA
kZit+TVEM+HckUvDA7Lx2w4dJ5fkrxcCzEHN8XocYHWHDlB7ZPQkhTp6QaXuJQGrx7BdClMQ/zHQ
WytlhkVZAhSUdB/yU6vCvDx1cOogxYuhnMObptGJQIQuMev2dEGPha+qh2rTn7vo1ho7lvV+5ajr
7+yWFBNd+rqHZfreh53vTEyAiN0/HSg+n51wtwFy9E5wkSzEO9GlyqfjrIdLzzm8yqCPDlgGZD84
bm0fP+O85UeTFkWPoghVWG0HrVpAM1uMi5L/5Tm2iHHdwXB9YcJehp9tF6HKW2QTKWRk30lNqcd5
6sFERZyTKRtF5ap0Yki6sJVPqebZkz2ERzKsvfunN7x2BuDGkrA85aHcYUMQvHAsvZc7IATQ7IdW
vxe5rtWXhd4KBYZctfVvorC2mzi6vOKq7gQqfWvYi8ohdHVYWhsfccPzVijCNG5IFcTB9RCWIlfE
wHl30TLE1GkHdEXBqVyxycPkeRnnSDtAwTbuI59l66z4iez24UIT3NAsCAVnw9WfG95sFMeenavH
B2/RsTf41ZHEMNsQ5Do9Y4xOq4+ol8xrS4J2N4jpixETbK3fFDKP5wDnGr8YqtjI/MimraAmxmsr
nBVgsuBMtzcHrq6Akk+fjz2QhoIY7vVLWb47d3c6oTiK2Op+Uqg2Kdsr8MfB56M+kr0kKTw5GgSh
Yt4oA07Pyc/yA5cBARddARNSlYietc8niVMmXbr8qWeZOOwWxLULueWhg8/H32/xRJdzytmDG2/Y
99vTMwou8tdzS1EyPjmWEaZurxTrsDDE/m1gqaqVTHZ+NQRzienhEYcv4Poa0U1DuLNDAjtZf3+f
H1IyQJVK1WDwrKJD/kcHOQ/HH0KupyvVmOhhp56DWG1iiOixZ52Cqlh3AUr++DvStsIe4WwNB2Ze
84VANyREphprOn3zaGbztNDkwP500n+Fd8GY2LiQHQmtyyOywNdVmPeOte2lGlwTHd0Wn8j94Aec
LWgYkwe5DyPAXbJTjIMaF7JztJOEN0VnkafYss9gfKjVG+2uMtx4y3P3EG2u7BMFYrcVei6MLM7H
dpKYpBYhR90k6dXQcp3q9u2isD65eGi+zlBEY7QwIO6SizxodRGml8phDHsdlbnHgUn1DhgHoUef
2Aak+FjnOxGWWGGj6+gUh1lXFSBm/UkL3wSeEGuuvG/RWyl5Plaqr7JvvWNsEbGezASOEILXK319
E/iVXU1XKt6glck2b9+cr0gDfdAPlY9QUPcjn1Fhn/5ZXHDquUNbi6hONFruGTvp+x/EB6omFoRT
Y8D4ZRQAUF3cyeK50NJ8hHuaz4pVgxXcdU2UaJQ+KK0OM14c/9W0gsWv6q203hLMY7XTqCdeqZm/
77kIIpgujqWZhnHnZNn6gbqPzZ8CHQvYSanLnWsf64U+/EnRlurwYJYzc6yse0X1NkwgwHtEdvS2
gXDO0PJCCtUYBxTDjmpJ3zO/zN/BarL89fcNGXHLaU9PO9GpntHXaepOLd3PR1e1Baf0Iy7LzN6y
+Yudzukwsc3Xl6l9g62VN29lnWKXDWzsLFv/LjWGzL7S7p1hx79Voo8GuUBc3FSUuGJ9MYtht9HM
RjMw1I7I5MDsqHy6jyhMQ223b4z0kmbU+2R0kc39XWMbcZSmAktEanDd3GH1ro21YdchevDfmTDz
3VQHok5zzy2RLBHInjtCj0yjeEi5VfQcaao+PUSBf91GfS5zfadN8XgCwV1I4S0QTPm0AnaHmDtk
GRj6n5qv3LUSiFhTFUF6la3c2vsW8vQ621AE99sSAdX0ibXapBwio+z8W22aaanhnRKSgfApovvz
GvBF2VzfvizrCWvvdQNXTM8JVJ2cOMAidrQN+wwnsKDPLJbaWeWB/GdY+ihV0H5HUW1j4yKUC1l1
sFySMiEAZVG+9/FTv3nyASXjAqwlucRnHufWLdL0PdKRYnAGHKaR8z4icbjdDfHAnA5AzagG58qs
pp/dfLNL5rAEcj9X+JTzxoOQghGHwe0YNooGEmfan6HGOOjFdULh8+g7n2+UmC8y1mZI5AinSJJq
bFHh0fJYkfWcr6ioZMY8TF9kztidBxcu9TkjA/5fcwxBCRWejAaxToLIFfPmMkIvVa6q5zaU9R4c
KFRp6BYP5eT1vx98bEZo/ue1zXaDtS73CASCzrgEfYaoEpUkBw+6nrYYb3h6Mki2GXcUwv1kusyd
0w3GtAuIzCiZjhNGI23OUcoEjJretEYlbkaowLldNrxNrzaPaAECR3Jo2RcIsW11bGqJEWmg7PuL
AlaV15DnIIQnrDZqUh17vUzaQPY8w4Pq9H1rM5Yu5xzEAgskNcT1WzeT1pXJgQfpZ1+Pu/3Qe5kv
qCGQAxPMXsJlCxxBIWj8K3XxuCTbGCdRTIdyj+Ak08f2fgNI1KHFtRglq8zpIpnkWuLQoaUha4I5
BHyQV0Zj+weDvqJwfpWaAZvM8YAC+mVMdrW3hkR0BF6WuwgcKwsRAaYg3Vvi/KiPuZ6ikCecDSu+
aajzivNZXk6qXaKblu/lf9r3xE4+IF4IA0OJv+BPUHZIusNz5MVlP+U9SHpX6Ww4FFYKr1GO4vrI
JPjMDdDN+/SiJ19PXN0rheGQ5gQUyfxztGsj4onYtAkqstm2iJ5PF2YHh/H9nlahHi+s0jPhEKXw
J0daCXg4LMtnF1208FMUcOq1psqOzp41VcJJEAQBz0n6LqDHx2BnecOrm8nyC8L2z4aqA/M5jO8T
33NlEfBTsEj0i63KbmQdxSqL+0Icrm3R2tEITTPU8AOuXipbapHL4SmgMs71OUNucyav60/OEzWF
bZQdbyGotoGoWA7Eo7UwLXyA9oA6fqjtxjtcR81oqMo0OyngJkIqshYPPcO98n5JDKu9sC2JmxpT
5XB7XC1vdSFmW9ke0ht/1lymQbHPhK/NPGm4H9SxoPx5WsuT3R+1nH0YSRqFiYg5gFGwyXNq6q4o
ySCLwuAekU6AOIwaejgFegs+hCXG8DV6DwUyKEfzkFnghRFZ2JvEZexQjIXXzQWO5kTPR/e7Bczj
kDv+XACzSlqTpNRPnqzpVa1HajgQcVLlguPVKhR8NeocJvHpCkd6X7VUVD4TZMnnjmk0MrK/t5w/
vH58QPhOJJERl+xkLTXiu+lGohXfY1fMynVy4w1f9MdsE43zQFE39Ss/0EfTGhR4AGZF5IHt3BM0
K9SdKGH+mdLPhjxu6BmOOLcNXjqdWa5HH+Rzx4UHVD254nDARut2sDQ7XfVmCoWYdanKw3coiD/J
eyMnWH41piIfKlYV5SAEGi+hzqFnLByaBuTx6a0XXThUU1QHc1C/NPGS7u3qt9qIxHJerfnpVz0m
pI1xRt227MOHBYXeDxs6ofU6Wk+jkASMJxzv5F7K+IHDP4LxqmJvq4NSPJK0pWAh13PbEQn3pEuE
SpIeURGccGFNxbAvQVtbgQ+XWuKJsjaPW7nt+Fg/X/2GH/W1H6dLrpAgSTkFPhSdXeFGn/W9o/17
2YM+yvdkktLET5XSrfaVTkYvE7glqfYC5Nr57NFVpuAPzkq4byLqJae3fkSyUy8ES9JLB4qRvocK
LCT5VDIydV3Q0OGo62eeliU8C6CA1H3B6P5X7hOgTqM60NWv+Crwe0mNHamgN8PykhgqvpZC3owG
CqPC0MjLwYNuHJQ1IBKpcAe8FHv408kR7KN4UU+XQUBN8m7DayYiXP2RKVAxeAm163Ylg+DwutQv
REvTKUcUV2RwebYAAix45G+UDkJHC18m5lWAw90ODV/ap4fhrZl3NTlR3t6LofCktxAvbK9QgiVr
Sy4TZG1LqBAJcdwT5zOnrArfzM7lT3NaFfUKTHT+mu/+3AQ1Omusb7qOZh36jOzK2jSlnZ2OD8SF
OyHDJPrFvAOl4AhbW3niZ8gjUV4qO4g9QF05hJa2AiuArrpSwTH7VrafXNokhBwMizyQa9oAHfsj
wF0VL57ljNAPuSGASc4iXyen7lV42TmzE4sfqb91AyN2G5F7NdbizENBL4fu3hk08HMXmEUkmQbP
IamJGObGcWizRkao2cZ8wUlsUQhRzatewdK+a7BKNHSIvGqiLzYNHGq8Z1NY++3I1UcOn1GLIZPq
lpoxsRRyPKHImuVPB0p79e1+BCRAf861uRy2hpLi472q9XhCewdweA9K9pT+R+Y5tp1Ij/Dck5D9
bMYGIGhSmUfU/n6mpJbtaePfMaxJ0UJnU6whCcnaV60zRC6ojoBtGw8pT9JuXFbGmSx0IU3PexQl
+gS9Dk4jtZiAiaGB5Bk5KRYGpYoCIRrWL/SdWcYZyYeXltTQU0gLc13dwPWw2C6X7S6Ahbq1jslj
KLqT7ndlMelEzeMY6I4SCskAZdYIRgbWOBFNEg9Kph4se12A/se2oZUYpU9i8gvLmXW6+cITZGOW
5NaVOrk9G19ZvinmReavyBVr6yGHX7UhDDkzl/p/CdA2fcERhNuHgtw2fqlMR/RBez9/dnLzOpoJ
21Qtp9RrhRfOBJ6w4Qc3kvKgIzEZN3MjWSjIRaOIm9AuxprLNdptNi30Pt+kH3qiHdh0d1+54efV
ihEoPxDcsCe15Z4qQYBnCcioBHxBwRk63BN/k2Dcmc9GcSsB33+UjUdvCtzYacEm3hS+pYsRnB6R
TmxfUR5ZCnlDFHKaqXVlEAEWkEMooZfyoGcZ5o8YdbjTaun+Ql1qFYS6ivPy89DtlqHNRCfwH/t6
G2XHYC0ksf0o42DuOXdc+2CVIfprEvo0up8h0mwA/XizWQ7o5iQUzcPvDSDdb/vGtIh6WNmybHKH
6LDtlM+cEl3wL+B7bOgAC/LmE2x20lraFRgKYLGEPrZSfGPftdn/Wjtkl9IiYYWsqDetcPWi6wrL
U79VD9K1dFP8R/UnorCz/URUi4uaLe9SRq/r91UKZGLavrBB15ScihUyYvscrl85qIYrrS/rEC0X
7O3/pOruRrbyW1Qsd8y2MDFe8PFRpcjQWc4xlsh5iCHgWo/5cUsEriBBmj+kz3BYZ1z11ASkkNbm
ScaUqrq0fv3NFz+Z/2kv0cPdaX0yPFM5J0npB8D8pzygYgW/V9HuVxal1t4bjTfCCoHELz7BwSbl
RVi+/pekjA1GZ9msAH4mamncVlypaFqklbv9P6U86PhZ/joeCC0uw26ORePV0suWeUSPi3Mp/g2N
yLM5q/aAKX5rnCxEmyJEPmv0OVVAHZ8nEzabRzZhdMOaKy797WJ23AywBQwIk9kADA3HFiZ2iVlN
zYGvDs9ObC8UFirbQljLLCFITLuOcmxxgZJ5Ieeyieig0wWg0Ms7YB2Cc3oVXYm2j2upHFpUhrbw
fEyajrBhPkNXVCkw+AzG8An/iKZafrBuYw5g8HQgjH3b0MwDDKvCdA3PHd/uinhuM0aOX5SjFSsS
OA8yJlBpd0NvTJvRY+CMT+y6k0i/DcwRCwtCSsfa9RT83QX/7yJ+L2Iirmxf+0pClg5+dSFdx9BM
Z4W7zBUIWGYlomavygwUpIKtZed1WTSez11ZCeMg7ldyKnBxzbpWdjrrIXu/Me+LJ/sTHKHrMU5h
5bkxPUiptMRXAu72KuP0LUK067iHnyzKq/L89Llw44Ic0SNnlovloBKuwcBN1L17pKT4X6AxcFaf
UofNwA3HvhF1lC27hqbPfqED9w2NSqeT9Lr2msukt5JzKLjYmrhbihIHvBqY21UP7rz2DbZfdJf7
f3HGnxaZYtScqaEmLFvmdBWGIJwn0CS72D1JYXdwP5BAzkfPRjmOtd2XksyS3WE17LpGdoWMOJ/P
atyX58SJDQP5eb9OSbG6X1CplDOXIUGZ0AY7Flzbb/rm+7zJfSR2iSQyfCT4QKGcP22DXnlK54GS
1zwoVak/3hYrItsLAuzvc63yoNm8cFOhg31VcR6KAXXNvVWEMDpf5oNV2gmguvwRE2cCCmBrul6e
/kQ5ymfuURtGHxv6zGiaETfn5fY2rk4YzYUWDL8r8o1dAxsFlO/nU6ZhUjo55TenAfNhn8tW7RYX
9HT2467LcRoSCBbmVVnUrs80BJcPS1RFIDgsQ0tW0wWya4QvqbgtszsB1nq/HKzMVn5a6b+calDG
23m67LuYy6dg3V/ED+MmKbJ8H7vA6sRBxMYrzT4TPTkWVTQmE/IMxm991dWkFS666qA9Zh9+NCne
RGsC24eFMWu1HVhY0mVCj8BRFQJZh35DGALP+zhEuj33ivenqhB+0GOJfRSo/3558ZiCSki6iu64
Kkwm9ywWyVi7ky3E/1OnIh8zUfNeH25XC5ysopHfquoO/Oq647lDFIr6k+kjHzjJWFIxQMmdnZui
hZo8DpQiQX0C5QsbFGkUaq4xrN0MrrOBqLQDuo/EUeDM/V6AQEEod6K/AczQR8wlKDYCtYwcoV7n
eEUE+MUO7YepmXblyDoVAqCgHGrwSTEzvbkqnXzRXW2aiyPRXmjvS26lO6y9Pv2EfSZ7NSxY3gcv
E2/HCDjz+mA2R8SE8UU2Vws1jfKvGMwGRShfrjdcCE2iuzqvJRrTtLN7HAbaq1evnJnJEjdBYpKT
UYh7NCA4orZDk4L2vuEwJtUZNGTfOB8e/DoxBfRHpZGVBCu/tfIE/DswfIJ5mZG/rCFwb2TZ6dR9
dKNMWWkXbVzwM9/IK4du3QvMfzC7SiXzMNxkZU9lPea1Lru5/TiagRFZPnmJan3ehHSSj5VAtBdJ
LY6SEYU3/p3I3LoQHRmFZ1sX6k5G8k0YOJqfUeJL4ERjWsw/GEVuku9lr0zPoWNr5jTAYSwNiobT
2FDidSsQ2+JOUQeMdxwFaMFjxx6xCShptM52ELd2OhBZ2tPQCdG3psmfuW/N87naQSxlmeSDcq/9
mQ9Fw+q2vArrF75QJvsCEd2uZyVsWxGcwRwHa/I5VKbo4fj4dhJJWs+Bu7yijuEZlb93PjXSicHC
oc/QXmEUxdaMH+e/eaOmssKIdeE95esoWyaozUqrMnATvt4MjmzWSK6khpHSrwZyKb5bl83iDQNT
WzdaovcpH5tEavClZCOJZem/mrilyvWmNWHmsKB1JO6bsgOjFvS23umIgYw9NGlk754oYiheRIcg
bp6lpWZ7uD1ud9MRJUzYfdUVmsYvcdh2khVYHE83HBIUM7fcL/gviLmPlZxzxL8NCGQf+fxu7b+R
cNaYNZtt2Bu15JAxZ+LIfj9bqhIJ9wPRF0TcilJGYOaGpHHg2sqqciA6t2vdKrKbe4CM0/d8agLc
mYbYem2zqxcR2XjYQzZeSf1A0BxPCd1a8SU/cj8gLNV6Lp/yiol35hMI7/6Ky5e5neRGzB78fDEF
A/3RfkMiIWa/Z9UP14sIFjtlemU7lWysAeUaSJF8ylhrgin/nXZpJUsYa7+OKtMhBpcUILGbWoTr
2spueFxlc0mzCHwG73beJw6Lajo8JOa5s6dUAvm7OguNBYRT/vTxgwPuCkbKBVPuZrnVQIcn0+mG
1MW+dOLVs7BrCk77ajgdJt/3gPcX3g58hCv4LMfJ0P4y8szD/9lihA8Tg2JRsHRdyE+tz6lG07Bx
n8dcCxGblCIyi5Rt1rbWRUwAijdb0ai6hkSl0ab6yHNfDhbQC25CYfiOvrIr26bXe7qfJmx9+KE5
xtQFO0xIu9fMbU6OgPKpbHg5GAjz4iK/2Hq6W/uUVCMBQQLm2zHHRF6vtKiPAwlLjZkR76BLpJN4
yqxrM4nfA81BfxoJiQ1ZCElRQV54OQUAGSsckuFSVfB+J3d/i8SVrwXqZw1OUebNAVsLYpoCx4TH
mBgUiyB9Yt+kxp6Xb6qd5Vhcs+USOqrESoXFhnBXF1E4qa6jEdDO9cX3g8ZPR36K8GO01Y/XSogS
60BdA0K9tSYHhdoqr+IDZ3PH/pVlCF9LDjN/jl9xqL9VPXPtQSf+AfqJLTz+7XCkGtoAICgMY6XQ
eUPOLYlkDPNF07Orj/Z61YGrmHdAlfsRK/N679LONEeHQyJVzTHH/X4D9jr0XvVbOKms1lamfC4H
Q8IFjvnGOm5drr/veC9U6YvyQco0mLsbxFKQvKYo7pOfZKUSu5VhN9LQKfYTqWNVWgSBz2ttGGQe
PVS0G1gNT/ELz5MjspB+rk4x2aaMjT0enwonbqXLXE/0A9g0+7MoTXWVR3/Z9d8ffuY46gKDIWob
y0k6L7P+PZ+XmPup2WhkrhTiAV7lLkD+K8NjnY7Rf9EBMBJMfk0REW3xXyEm2KJdIq7bhSutpSAL
NOrqs+CguzRiNzgT2jeccYd7H84DxsQfWoJf81d6OvQhVO1u35tf8PkTFfYpwXyzzXyeDslYu2zV
/1byflPLJ0HsVsV2z635Llgw0Pg2fPwZUZfsW3lZM+ELtKch7/iG74/2syApJ0XRafIqUyRSZDMa
6Y5bc0sNFhiybdOyOVcDf2cA7W3N2GIS30UC66nNgdxwh1OhRK/Lkhpz+3HT5RntdK2RJTv9z5QK
fT/5uezjMnCKwpNzail5ikVMRx0PSuV+Y8QZLelb10WsJsrHf9uVZTcAJvEzDT0R6cpsTnjl/FgG
u/KW1cBqnXXxM/RKqjXEnhcCQpGPvJtZz9Tt+dychcpVyF2CVN1NpBTQ2ZFbWe3ZYWEtOQ+gObDa
bHrFYBd0cJ4uYsV2Q9wM9/SycDDwR8fIu3j43btkEE0xrvNWRlSgltl4DD0kyB/svI6WFll+WN91
kAZoVxcVJ9P0t50zg2Gr7NkOhusQp3aQA8/ooP37Sio5vfKBdDqARs6OOjfB16P+/924xTfbKqRw
/6SVn2fX8v5jwX0niFc608JtK5ZvOGGYe51gYVVFJWGQ8T9cNDIUzCOQLn2Ohu6hv/yzVCOQxfvv
PQCc1t00ExcLa6fvXU8//FBvR7AVWA0U4lKKi5sb1tPPSZBTsZm9owYqUcjXocHYGwn+QXdAztXd
wv7ClS62TYqb6CVHE3GIbyCApKymCnazcgzx7skQk11dKKu6lPSvdmOACBYqBLM3Az1exfaAjrk5
/Ps111obTG2dL25eR6m+emcqUauydXoAXOAPS0LfT/6bv/bzVhL5wWVvvwIi1ExUEEmczuBqWEZQ
sf+dAyJAxMmaWeivC3SYGIw2JKxiGJsP3ijD/l9CIIGgFruPR0C3gxG1ReIZV0IdgPEemPqer8y3
v1jm45WvYnCFJcb+sWa395wU2x79cYYcv0qa+qmCugE9dFdrpe5huvJQMnsbZLlxvP6sOzZAp6Gd
Qf+SSXaBD815EAn0zHIUKNzMQF3x2AsEBLMx/HajpOgV9x+GZJDe/bLj8fGSpTDaGhy8aSosBIts
cZxH3GyXhVNsDtm1IReJISKTgXPPM1myTmh1o7/0cEB8pNDQYiBxeYQlaKXTJrLRVDr+nfuz5cqk
jG8Hd9ozhguy20WOAaVtK8vHDcYLjHwubeRmLwYjHZ6UjKq+224DQm55PqCrKLjW8tBWGV+IUHN4
8GSjIkTBvWH0dTC0qqauOnadyTH4iN3vzuZYmUZkaCJr0SS4HxUysAXGXL9f3jJUXmW5T6x43ilh
j/ixhTSTU8/KH4V4ANW7+cZUKtAm6wFW8b+coj4UlVNC/QeSW+xR+0dT6WMsC4InuB/aSVqKgglY
tqJeXsvV2VOmi1mRc+u4UXnZcf/6EwXDcGQJmDGY+hCKQOb3wjsmuoKQJ9ANKA9rVuayQ9lHoukA
MQEVhIk+whHCL2x4KQNG8RWp1ODPuHFLneoBpUZ7M5FC++cyanBR9rOddyNZe1uwaTiZJLBxIEan
MCj/03EqbLOGV0VRp+w4OP4NcuanLG7pgurtJ5DqhV2fEnbFNSL1PgGUsqnlRzTwNNHdqzI0QV00
S8Sh5QZHbsiLf5czSM1QXaIabIDKFMbDQiCLpJ+TTXzAeRofQEk1xUUhSWrP1oifquLUMIiTVOA9
CkDWr3D8c+KFG5kiOsP29vadYos+AxRo7XObN1YAAbg+zry7w/qkgEZcDCKtZkITt7OOawVyoqju
PYCXv93AYZqK/u0izsaT4Gfq4CO044KN/+FF6CGqd3/1HXOrxu1lEOo+vAR0CIHZh/I+LucIhXdb
Xl3+oUQRDUyRwnRn18NHQPRGcSHUT5fYeHkcAbSeyB3FIpKcJtg+O9xy/Kg4hkUGeBsLxMEeUq4e
iGlihKA7uJstcXqXDYVw/4tyUuJ++su6Udz7MA0f7mB6v+8jnFLl/WLHOm4v6gCkFATuvQk4cw24
w+gMtjWfWdvvkOe5lFKU1n4e+0aYTWBRpoT0xpffsUp6nomSN38L/oBaqaLqiM1I8nyjht6Btv+x
95rIkrWPS9KL8hNLIqUmIzP6BAFNKEqKUn9ALmNwwz0DA22ksDQdbijDyQE9M2sL3RwMqVbNFKxC
bwfclEjej7rVmVLWEd9lKGVpicQzsaVF4QTdkvZ3pWS+A+HV782aZa5AjZMr166ctKHj7/zL7MQZ
mbuXi02B5AWkXt6RIV4/4bXEOGZ9ZwrfARpG5vVAvr85Pq5SiR2723Gmg14J9USK85Fnb36ge0oZ
D+U5qrzCOB67MSZemZiDMIEvGkYu7YpHWy712hCxN8t5spsx5QYZH4kXiRayDubnO09L6aTLU2Nm
fy9k7c11PQdIZ43y8+9MdoBMHlXxW+Bhj3PFHUhobUfW2WFR1folXECx+RZuFKrmaA+opMiqYoDL
NMLzbzYipa1hvFBgljiC73iKQa5ncF/PTkgZsmyAYaM9yBRfwSMRFQv8lKpYgoMYoLGhZzkmy/tV
7XpPAZTZShdaK3Rt2yWZueKS4mmR69aeGGDtAPn8EGVa7dz/UWkbE/gGypfeelzJ8BaC6HyNT1Yx
BldWJqXHFY6upPoSY1Xleod/nvienr9Eew46fVNwrsLTOuFdOqzttkuuF19auMEj77euxmhQxbS9
EJM9WSDDhKl3dKssdq+TeNv1TADG8RKzvQn7Hk91Mso6ztt54XyVZD793i1hyb8fcWcdLJzrjesp
XRI6pTFR3lT0j3+de4+lJT4gI5GrQwX33XSvxDoXc4e5+WG0H5RK7OdmfkVN3Jqfyt5BpjkrUqmI
F8sh/1+gnkCLzgctww2CHGtcO6NfVEdDJ4I9ssnrOTAegeaTMAcc99mBJmdwNPqyhjrQfGf06GYJ
WsbkS8vZUUnF2XTvsjEfTp2yg7JxUSrmVsW9YG6L+AFgzVJhJEHvXTHLiK7cZWVkQSHSY0Uug2wj
Efe971gVD5+yywCU7aTRBf+9bpuI4ud/vOmdmrjbm/O6XUrL7WxOXD+6z8/uMRrccJskSo6vbO3M
QovBSsqzfYwmWpn89OjrusBXTd78q9+mMWkIUO4lPt0ibJBmKSVka4XQ5tkhruopdMWvfDAjGLH1
bYxYcwGfqNLId6ZJI+/xgDsG4kBTh4ApniEneRC5PusVJ8NsskPwZ9TRLCRJAY/yAVuWeS+W1h4o
N8cUqRzN6+4hmgFn9z+kR2MMGGhVQFc2FUTqRK/0p8FXxo89hxVRIeOtA4d7fgrUYlV35LToBzKN
CLBG8A/n35R3OCI5cPYji185hE8dDo6yQNfIsGNXVsuOv7Ep9a6dIWcv6n1ogwPlKCCgpwfmP5iE
Y3OW0Tb/now1oeT4pY+iXVAWMEc7Uul5aU8SP2CmN++2eVkoTI5lPDKApFZa1Uk9brkLh7RvV/3y
qfoEFWQiSnimIveTImgV3Qn9ug6f3I8cdqianPfcrRvz6iiQwYFmUq643EhYH5BaWO0NWIEiueEf
M9QUAmfyhhrSCj4/z9fdvFamc9dgtKT5V3FaVYuql90Zf4GPEWvYgitCaVcoYeXSY4GYZZi887rz
mdZJ8GdMGm5uyAzQj60qpYNz6E12SZXSR4XOzBbFrEL9U7Yhs8A6OlL5VMfg7PT0GZDevCvuj1ZU
/b33VWcNUgn1jB8fUFMQvwnvxfc2RQpn4ygHTuE2wOcmlZmognrZ6Xzl27/J7VGI80gwjWjvzv42
a8461h+ZZh+/qDMSQk0lj0gHQbXMiYGuwCCWMAbT55pH6q+95jLdH2tZT7/ifOOgc4EriLmriv0b
59D/tBZTVK5SaLiVzgRu3VasR1hTAChg0G0/UDnIIiWo1lZaPYAoti15btz1uTzEvKNgRcJxmwn6
czhTJbga+hEew7S990FCT3NdOdsvJqmge/hhJtwc+C+dadf+nCSDjdp57E3P1ZvnUQNWfxRdfHjT
u3MBKpfk6R3NsLtuvcYkjeag/ZyuySpS593i446V4iA3Gy1bu16kG7Ture82I3uJuNubUvVTzkr9
BGodMd5ACZL31IXPoDgas95epDUDLZWNWpdvn9b2+G/FyhXNwidQx3uKoZ373obbrLoBItfJ+K1I
SFJ8JKWpKE6xOVJcM9sLhQAa8anoGt8DLedXl/SnBz/gDvbcFII3flVwfE0qtsThWdbt5K1+2+Nj
XdmVooGgEC/9y+in1vZNaB5YUlsqNOTOsg2Hmfn7a/NDpCsIBTj25kwPIo5a08cWeA8qhJpx/cdO
fkeE3ib1XoEQXiit8OiTkDN0Anyx6bQOAHgRA5hY/iZh5Q5GrdLLeE35Ph9nGb+C7J7ZuIThbpdm
6ePnYcRKDiVXKI+f+BXMFx9Yeiykjm/7yylPKq9TsBJyEgITi4xEZ0NuTzLS0o2zMBFxD035ffi5
dr74OXCLlZQfZ+2gTAUMsJ9gdpUMt4QZtBJFePrkVjYMFGgU0hV5ISRGx68Q14f+JILgRw2E5r4w
86iue7wp0oNjCZdkH8Wr2j7QoMp9W1zCt7RKE8fkyRl66ghuSg+vOiY4j+6Hp+tv5ApnjlskBm2U
VAENVSAapQsHbHaRPMUrGJTvrRD5d+Ses+kcbHewK3pGYXbJvotUj6waTExUY3Eqnqho5mofsZbT
yZNHCvq5M1naMPamMCLlRsnHD8qBWAiNjGLtxg==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity fifo_256x512_16x8192 is
port(
  Data :  in std_logic_vector(255 downto 0);
  Reset :  in std_logic;
  WrClk :  in std_logic;
  RdClk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Wnum :  out std_logic_vector(9 downto 0);
  Rnum :  out std_logic_vector(13 downto 0);
  Almost_Full :  out std_logic;
  Q :  out std_logic_vector(15 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end fifo_256x512_16x8192;
architecture beh of fifo_256x512_16x8192 is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo.fifo_256x512_16x8192\
port(
  GND_0: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  RdClk: in std_logic;
  WrClk: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(255 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Almost_Full: out std_logic;
  Q : out std_logic_vector(15 downto 0);
  Wnum : out std_logic_vector(9 downto 0);
  Rnum : out std_logic_vector(13 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_inst: \~fifo.fifo_256x512_16x8192\
port map(
  GND_0 => GND_0,
  Reset => Reset,
  VCC_0 => VCC_0,
  RdClk => RdClk,
  WrClk => WrClk,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(255 downto 0) => Data(255 downto 0),
  Empty => NN,
  Full => NN_0,
  Almost_Full => Almost_Full,
  Q(15 downto 0) => Q(15 downto 0),
  Wnum(9 downto 0) => Wnum(9 downto 0),
  Rnum(13 downto 0) => Rnum(13 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
