--
--Written by GowinSynthesis
--Tool Version "V1.9.12 (64-bit)"
--Sat Nov  1 17:22:57 2025

--Source file index table:
--file0 "\D:/FPGA/03-outsourced proj/05-panoramic_camera/cam2dvi_no_buffer/src/fifo_top/temp/FIFO/fifo_define.v"
--file1 "\D:/FPGA/03-outsourced proj/05-panoramic_camera/cam2dvi_no_buffer/src/fifo_top/temp/FIFO/fifo_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FIFO/data/edc.v"
--file3 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FIFO/data/fifo.v"
--file4 "\C:/Gowin/Gowin_V1.9.12_x64/IDE/ipcore/FIFO/data/fifo_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
qEoXywdsfxwMCzzvkiioDdmPGA63hmez9kGQW1+JwqsxKPt4zC1OAm+lKnc7b+JhQMWr4phmlmd6
83GJyqGmQRN7omfuelOQ6NRha2NSrm4N/m2fC16JdJoqz+NQb9CBcBa67SrvNP/ALLGRWoyowL6K
b8/5Qu1+PFGnIwXOosVMf83qWoDG6Jr0G7EJeLTI7/u7ZxgZHerJVuav9itZhM298ISfv46jO/7O
Amfe7rAanlUobnAZolWN7/NuU38v2w5+Vt/kApQ7DSNTnFwOi7Oe49YX6P8QABKRTriWtDgsVvn/
LsqccWC17ZymmHK7MaI3FgQOcx9/gnLLLABLZQ==

`protect encoding=(enctype="base64", line_length=76, bytes=50848)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
BbXLhww7pvAiRt93NV3xfTbisRWDNVBBzSbOLmaw1XkhjYzsXB2brlJ1uH2ekXDKtvi8IxehBWqp
Er77XJQ8MJQSUSWnNBZr3B6KxMPgFqC5ZCcbW4iv/q7zD7C07Hz/aE0/P37qFPCKVGcn5Z4Lr1S9
257pfaAfe7ZEL5Ytf6cT+ZjVMjQ6u1IxbaEAh7abvwkLbfAZDZG6ne2DaP0yAddjOIvPNMhVEP5u
P6Ljz0F6xx48d8gnqfk1GKNgOtfLgnVrdhiv4G/+amnviplqN4/I0oBRw90R3mbZPvvjQjTceUUA
87Y4Ijbza5TzyJ1k1whGtmSe9L0QQYCyyUfsDzi09KJyZ8OuzIPYV6Y2iu70cAdXau5sLlWZ8atk
UFURaer1vAGdoFP2TPr+xerVhxyPyHMc9CEGZhd/8hrqIiX7nZT31cZxZM2oH3kzUs/TqIJqnwq7
bnM4y0CDrvHcNp50WearrgO9wNb0VSvR+zCkYgkxCZUHKA8AVOIUY5U/9Hj7SwkZU5A3ubrK+Cjm
F47kGQ6l2gpa5mcsKkGGOYlPAHlWpZ5Fr28mjaYc2OsPLUpqKtvHuU/6c59tgCcBAE5fUgdqgzEI
Xfdn/QvBmuBIoZLRO1buft/JBDt9kqNZ/nOCTPjAEdaV499ZYcxRBlA0Q4jdKWo2UohhV/SttqtS
R6sfl3J9cshNiYHW7FuExGNb+poyHXBzCz1/ttY57zGVQqtty/nShDvadRHL9RjEu5EWzMW2sPHu
Q6PbqDrYw9MbUBK6PyNUT4vxY8UKB2PnQm6/DxWveeWc4y3vADb0hbrOFMmScTu188xBralw4e6J
MoisBtmsgGZW9lH5EXeGJKyAdsOamIZUE2McV+brUFDa4430FbNrYXxOrHGy22Wgcora37kY3hBD
25odBqtvYkYtdNzQ7ysEr0zJtm5+XzRrOJycKhwOtkJ22nSgZo64z0z5j5UtloKE1MScRJVM5Maj
2dDtEUuqhBMmOaAmdIQeCNJs6F1+vyzNVNAyU4F6lcqu26njakpdRgDMfTFXQdhqlpaDAsPJDQXW
37GxKSB9jfAZkLSvdzMgSfC+mitqx3eqV8YimEcD9sXwGvLthuHEKwcNKm4n3GT3SeYDNVvrLzPz
khahpBz4RX0sFCPUYWvvKhBSOoYUeWomjcvyDN8yTfszAFMIFiRXOXwu2WoEq02ga+TB1WZCqZvL
GKT8AmF/vq3GRr+WWnG4C7Eo7JeD5Zqhn0QU1Twq3HpmGjIDASBoxR79qCKF9LHIYkTSM9KWHl4u
UTeTVMXfzPXg7B5NLuBdS+yKUE6Dc2W/YoG6ZHnCdZ9r7b/iLMLJfX7ne62dAjMB72sbGec6DkAz
qTdFExMEsK2f2AXBr9yL924LUgaNsBMm/k7cqbikBYwdmfyAFBghn+NKZXLuJZTS3rW37MCfg3gv
uQzoHlxqZvKHZDSsU94SfiTpWNO8oJe+dWvoACHuvWQadrIRfocLne1YzmPFD28ZngKysOn9e22s
NYVi1JmuIbz9h/lEAsEuKfIk3nPb1RJsI7g4dp54u9M/kYwUNXzBhd5X8y2CwllbrA/RubJB6Kyz
vpHyzXhYWYL8L1DN3hZacvMPqKslNE3Q8c0CIQbYcVCYyEXNCUpU4C8S2s4+D3rMF6nWogyBaFwn
pqIe3XHsqjyS7kWy6b/Pr65oSrjbxtSnli7d1Oxxvl8wbWZbE1JfV3XN8R/KUM4QIwHOtSBx/J4C
PapCr3WhN5F+V5BCOd7zEROhBi6L5CSFgbn+6a1KTAe286fiS96xRYFr/JAowLlOZdjK8sSD3Van
InYZbdUzG3mCKJjnXaby1zyVgpIArZhXIKTyF3tONNj5OqBFjVrGJ/Pe9d3lDOChgKGy9oo7ymdT
Zld8NfMKoeZD5jiOqudbpLNaHivAqitdUS3AI0lfUBY488cFh9fGe1cijAOzZ6fZYOtqf+srTDZC
hD8LKlcDjLWg8YIDE+wIiAuX08JqPNp08ipYgrxWwoggR1rkD1qknlPz8z7QmeWLfzkNn3fM4heW
erLV8+gXK64/TQThDO9AvuXOFUd3Ntowna94AlZSF/SZpXEwn8QGpFO/nNnm5+23n0/OaDwPgoTj
9VmeLCAdl7/LscQyj7ySa5XD0hxF7xqIfQm0Wzg/FwlfsHmM0m0pbjEXbGJmXz84QlQYWo/2+h+T
i8SEZHqMZ8DS4cOR21QMvdJZ8H+8obovAl8XjGGL4qxNgeMAJUueS7ITHC2hoT104m4n0VR2XZ+Q
jrIJyOxvjspWysdqw8dEStycQpXZZzKVKypXTqEIrBtwrw4BQHRxLj2hcLD53sHbAl5lMNCqiWfi
DMR/UE2aOXqT0gMKek2wnSj8F5zBbiqRvlByMbzZ4ECEizxZF8o9yC5bCny4pkU3EV4OXGcDyx4t
lXRXrHB8V6592yKHL2HsNoG/R9pAt5CKupJnqLza8RyZRXj4FIf9TNIxi/dDjUeZANHeH3Y8S9Br
YzESl+/8xK37CfHUJoWlwbW1GDsDWy3w8JJCjrjPOoGX84F7VKDsSkc7Gomgqk+y2MiVKLLJNmai
Px3ZUqaPqCDZL/isCsr61z8YEvOtvThlarNYQaT54O9TsLnBuFy/VwABjWpRCCZivWqy58/EDBID
8xvzxViCNIAATxuKQr4XhQajFd1f9OT1S01l2xMcCqaXPSW+IZa2fsBTAbyeIqbRTzk+rDs0FOq2
yBvfu0Q9mQAhB0r1zn39Ztiz/LQwyJ8Pk0wMIsoEgrX8vIl97i2XH+VnSTK0daYy+5OxrSdndjBW
niTcyjyUu/WEUJqj/HluqJfr8BgfSPDbeEKSpf/QfTUFivGia5h2jCvqU7hWhmTpmCx+Kzak6EHT
FNAdW5G69HMK3Ihr673dXn7zExPnb9DmrazeHQssV6/0QNEif+qKh7fl9CFLsGBNWXtwBAoYwM/y
f/nWJuibkYhCznNAt+LdZAWu5B9Uh1JcIIsyU4+UwFI7GMvOSKLeMB5EHDbAb8Z/hIeafFUdPca0
+BioFOZyfJBAP+QADrZgahhbabIFPJQOUcbb6FJm6cRTmNboejdTgj0Gkccgbs+szWDlQk2RaFHq
x7fLZwbRjoKLF/LtVKAHoOWaAlAPtBH2QI3eDwBwgRN2Y/nsYGNp75Nc+v3uqKsDBvPBghIk6l0q
kw+V+0o8ixth9YfGls/xCbW0vNivFedu4oETq+k3DYjfk9d0q1xAxELqYsHjfrOtxKZjHZBho49G
eY8V6fLvobLXW92XuuX99lyY5OJgp6/ghO3aForEK+VZ34h73HRKQqZYPejO3fZ3GrSveClHMXrv
GafLx++rS7JteK094PpumZJtL2thm/s0M7N/kxMlGuX7YBo0ovh4QFxHK0U0Nz7iHT0Y6ovgtP7a
jp+J2zDA1HhHamAs6lqsLWpmMMLPOdi0QtMSDY28+KlgDKfYqpPwic9HWVw/k8UKFFOOZDNNi1Yl
C6la14MpyeQQ1NNWH7ZV7XN7RvhmNgGcsdVHRjyH8D5P/AY3dqeldExQmCc6tMWem6x+teEy6KMI
d6fQ+bzijuAoY2103+rUIUopn2+P7eSUKW8MPIoRORj023s0pWj6rp87QhqYaLDlPhenvwBSIqfj
YYOWecjIFnSlKwiqazTJDNE4BiGZPIY/hG8aH9Ciy+kJWOq+jxEgi60SMsW75vERjifIf3aIO1XB
9gWk7VRSskO7zRpDeitB2rzvpm2KiFLd5E46LnjlATArwz54ujq2aRH9m8c5VYWkwIto/aaJoljS
TPTIpdyxj9zVG8PN0VnGkevwTxlyDedq9XgKOZsx//lUBOVqqRJxu8khfrUNgydd1oMzx+/HP6i5
XJ8o7IuOt383pHu1ARH75Iq9JTWzrzZxQOdiTN6nj3Z8RCNPLI+TNp5GvYfycxw8cJ+oWZrXaqp8
oV5iGbOVXqz3cV6Ci5i89p+CfYAgoVnUe7WU2sxYu/9SAqzsg6HAtbEnrJl9f0pGLtSCT40ihI7S
qeMIDevWNHBkXsKozZZbymcjzPnhtxRKToPFxtv9Q5cFPoILlViuOaZF2gmDMiTw8fYwu15JbSrM
WoLx39RfqXRGiBD8yKfE4sP9eLaOfbsHXqLe5Rk1TBGbmGxMA2PIu4FmnM2f1w0a5XyF+821BAzQ
8KbApDM/uMzc+nVY4ptbcNNi/EuUCnB/pdNE0pd17SbsXf02zm8G2SE7LWih3xi2+AtBa3G95RXy
gO27rpH/8JXJTUasO1v+LFQN0Sd9smGJ1PUeAEaX8pMF6vJ3IQthSiNSQox/6LCW84vMu9LufvQO
HiqWrmGNEGEHimofLE4PoEpnvjSLaCTxNmKL9L7rocCaEBv4yxxvpaq2Ufvl/nxmw1kg37TbJ6P3
GJR0jLTMHtiWHkhxi15j4olptYRjdAfocY6qvzjiTv9bHnIxcWkB6UCxC81Hkh9080Kux1l6E9Ch
0o+QrTIVWbsYmPaNwfkgdEauJdHZrcXyPUTZm5ZjwtEoqA1kI7AW8t01yl3am2T7GLVa1UD090fY
ojKGOJ+pjzYQwnzhuZWU818VZEil5IDHmnS4p2aHGiOyyoDn8AJEo7ebFTuU3KhAwONBeLPuZwUm
G4vNJTTI8x6a/dAG323/B9D9Tzm4vjZwZW+ZKzbP1PZQBVXCh7T/V9lz4YLP6NgB77PTbT4hOw0+
c0vumtJx5fNdnECfgI/FicDG1anTFo4ea0yhubV0KvanX0kaeTc63r8s58JxAPOpJy9kVDQmbYqH
7YFjUEmWIWRwHe/vfQPjtcqmuvo896iz5b4ToIWwHv9QdnmEzZXyw/+RyorHiYC/87qDboC1zUUq
NKDbaeEvbCo2yz+q5KakdkDmVPf8U7d9Kc4atYUJ26AzE1JMuyKi+5u8J+fSXFtt9CVwbpGxcrrW
Bz/TBjBiHaRbXMeGF5X+J+CH2A01uNum1Ov54C44NGjnUgomoiQfDv0UAOuIJHQz5CcVFWArKyuS
cMoEYENDpxUnrOT0SWlpA2YFq3INRMuHt297ugXNPLj/L3u7ayq+eeq5y1no4V3vjcUW51wNUb1S
oHG16s1dItzznMm+a09Nee05Wf5lPyXpihwrMBX6vi6ZIX6mCoaOwkkH33DKPuAbnAdP0ghrPY4s
5+GXguJx3A4XWLobxMrUcDC0Sr/0rDAExDd15UCraCfs9e/ngR9brZEcbK+Cx7FGdI/bkyU68igZ
q0gehjtOzgwOf9Th9i6ieTWjNokSQXiksxxbNSMIQi2hbbyhS8hEa/CXuZwgPVVWi1vyYSR3FKsZ
2tfhKdoi19JbjRwNwvHmiSeIryqd9Pr8EhSk5zt4dWyiGkMaNl0dguAhl9vZBhFuSPqbbO0zWwkr
owldvSwETCbvyArxq9Ee2hxnpT3OA3rThy88C659jr8DLneAUJYTQOCBPbq8SjBBySkgeLO0Q5tp
GJCLcs+CitWOe5UYkJmSXcGhUIwc25NVxn3U9dKh67bsn1p7yBY+Xg4Ao8M5AgYmYOrE6Hj+EUj/
YgSVm25KZHj7stmqaK0SPuKtyppOTV8xjzZnaqW6WWuN8dCJttcD8sXb3yFp+fQs58R7gr0cmFmv
Wq8z0AJCS9/wwmtqXJbfyAN20cAOYBSqfF3m5yI+lgZ55njrMhxTpu4zoycpMg+mc2INvEKoRhGi
/J3MFoAQZo7FBJceFPKWOQDFtSHCRR4+n+OiuhnrXxv8pBlCLgjoCqvom3JkUlcUGqYd18SVu8wg
bqpo7qzTR1T6A+zasbb83GNOp1nsKM6w+ImI2ikWCpiAMa3BXCvTEEGDolscN+FC4fgD75ZP7XpO
kBYNxFFO18PgtkdongRvN3UTUZKGMh4dB1SCPhYLtUze/DAKpzc2rfssizWRKCMlKdxs0IjCT6xW
0smmODM5MiR4ZnC+h5XAJ+rvsIPUawmBaiOm+DcAAYIkOaAOhvFX4svM1jWoOHklin9/jNbx3/Z8
In9c/TEuLwkKcve3yGx/Pe30nZ5GAPXPuPDyaaQfk0il9/RAggHmJou2Ww3n1+gHXXPGP65BjPku
FJbUcPTiqb2OxiUP/VL3jWFKe7YAj2SVMGLiwLL2I5b+wyCHxm5Tutfotdvtn4Iw++hJflviBT2n
DGqVdBVZbCH8o/EbAmx4v45MK6RYfWZNd9MWgeHSOtyFlxh/cQ/BANdZDW7Nhy4pPe3hQEt2UxfL
Kj2LJ+DFyzp1V8Fki1hNA4Ih639lkSvAE/qicKRuehFzqbz6YTD5g9RuwPj/HRrAOwHPPFNmdNJf
LYpiSuy4v+lOOWnUrtI6WKgSv6IEyKyfv8vHnczHufcf+rx3Nsy7le3IPXahDGRQxjqWGKAGBCsL
Eo9CifU8To8T9zASqlNUG/mbUi3f9PqV3duoSnTQCbdmY8mhUiEGi7Pilvl0GhJvEk7OxvcMbV7n
hwrYCGgOBC1Hp8WFVjXielVC/pCL77WJYq49QjTxpZ7HUjUebjPcikRHhITmXWKl3klwn0NMtVuk
gsDDEJ83SiDC24Cc2E7mUcZJSXhrC7HdQshb4kPzLtFyZXMiLNM3SrdcKCxdQgO0rwfw52iB0jo3
HRsFAIrPthk9OvKdU7tePxlYSXXrx3UT47JjoZpWkF7Lp/5lk19ru3PsCMEVhG90tJQajMguJ6mR
u5/mBG29Xae9xZSpS34htBleiR91mRzxnh2ntDrwjW5WoOeqZtP5Z91X/gbgfERSrOYoIWWqkAUe
b+Y6Cf199QxfRq1liJ/2Isfjq02mLzcWjmc5ESdRjBKW1B5pw37uqCWw+E+t2CpvXuvtahSo/XZb
9PYkVv5PiTG8lyngwGQS7t8yIN2nvCY4iblqoVJj9FPFXNtd/EdjECasHd57kzLwzegcEQhQbEt+
ipxxWyt0dikHeSKNaULsXcX6w89FfdO00x/6wAnfaSCYXYIpOOJ+FvZN2mbobJdW+l15uYo0qz0S
hG0P2x4YRlIW8k5SLYpwiDK5JjIFTRdoQwnFRXNcrGvuLD9zrKxZFANi8s/KNtWDr44qt8x/F3Ws
kX8oqgxAyY0lqXWjQbSzK5MtzX6Wgh+tP1OjRn7XLFBb1FAG3LDHMAUnPyO/OLyFSkJxGgfdmWsu
q4qlVPfRgRkAaKosZ775qeR+sMy5xlHTr2mEkky/qs3z6HL6GOrjydq+8bEu7KYowBxK19tJkHqL
IlL0VPvfikV5B0Y7Pau1JgA/nhOI3BjKoyldE5y6EmjCTmvrZGZYyCiMdJx6q83CdGxUzHvI+XmK
UNk11x7nLPAiYI5ZF6LAN3PkSGESroB5PTDvCS8UzzRJcVhLS4AtEsMR2zhG4yxcLQP9Orc7siy3
V2AzPbrdgHVpvq+oHpIi7bJ2UneE/nTkOBCG+3rpszNOIiNs2W8zqdb0kkHO8ng68e/Ms0oLz6CY
HYaSWe70qf1kKKWfpZi8lWa1Rnw0s1EtT58LCFwLYDQ8kHEpywO/eohqc3dipkfQ59+qTtQCpdQm
3+NyVILD4yOWdzfZFIL/yuUEXUbKT9sKDzJUBMk75agFwhbHi2ir6gM3m5trzXYgm9BbRYSwdcQT
0Iby57B/BudZrG/U3U6uGbQ6eXfRzMVtuovxkoVdV0T5eONzjGXbu11q/7Rb2YCSWfZfNyVdH854
wi1eNsjtkvNSxtnicRNPSJ1H+VfXKTDOva0/eTXAUAHl+Br4IrvhGSUn33yfvBTstpXf4POkrCsy
y82NL43OmsHRtlCTQm3+bxIOFxUyMXMTsIFKzYht66luO2aJ6gpWy89wXeDi7r5MKYdO6HEaHsOU
s6fJJ+8il+k0LKMNgNvyp4euf7vZVLolzDo2OY3WLQh5SFti9k48Wz4Bi+2GIxMIUaDTMQDwNp5/
iCsaYRAU68Pu55Ydj2thoqyLb51mBdcvagrgC0og9IKdR0VmfhTFXH4lqAQ3Uuxa7LJ75SMKVXNJ
rBDYmF+6+fCZ6WXJfjphSqXIwgBdfIv77XFf1Gl5BGQD0IdFVeL/49zJGsIml3GZ1vd2Y2bOsyYN
iJXY/8PzkXOrhyZPfri+KnIvGVSDqUDZAE7WuHFrsNqs5uttkXLIOM1bQcyWlxdPrcmKMgDRQ/0P
7knmXwD1DL0RDHHFAueRIWpnA5fg0zGo3xTRuwHmJTpfVuXId310lT9q8C92OTMQFFplPP+l1jDV
srVOcnD2UV0dxRBd3YGX9+JfE6dpCeqFaug4yzirwlcjNTS4tXLFVE7KOVsZWU4yrhvQIADDOWR6
wwVEJmZH89eNxuHA8Qz4ToLLh57/7E7ievFovZBa9lqMZcctFGbr1PyFhXdQQtsEdOZ44rW7W6on
1sw89GmF8onNWb0VtULjiNgh7tTNny9x0VCcQKyxwOaWkE8cokbb3YhMiaoUpZl+PJv3u/HW/FvF
fxnxnO8An+A4OwYC8hOGL4jYumpAHlBzfeO8T67UkrR55bF21fuNE4Xvn4b99+YbTPlqguanryO3
Wnvsr05tKzjVLmvMePZ8SzskdL7kXYWl+Y5TqIsiU/4ZiuSBji+SsIoz2WaKYffnKCr7KsqHS1Fp
KvT69OI3WaiTYFvhL8e1ygdXNbnhK3nWu2Qewn/BWNc4UN1L4urJ81kyL+kfFHkp+5JrHpzb+p7Y
3D1L6nECsizi3KUYg7EV6vvhx7++uW8cVRRi5e2ubZL/evXrHZ6mA6Sq6mD7r//8SHiHdGxq6Z7Y
/ZFbPjcnSqaFL21r6e/vl/ptEF6s0bl4/imetyXK4dIfflm/OPIf+B/keQFI96rG+hWcReRSfAt7
xnp45zNYYZYtHv4l6EuvjCQxGNEAgZfMjU2BJYa4/uP9DP7GAQxw1SQvorQmzanHEuSoicQ1NeY+
9peb/eDDediFTNv92sykh5JxaclxI4BhHgLpExHuYOYUdxJV3gLPZWvhHa4JwAAbmsLlcMagV+Jk
7BKjbTweEl4g9BV+eBnN43xTZlmOqLZRZo2ucOHszJgHfnIVQAzkIoXT9/xW4mcyJiI93oUyvavL
cQ4zWRnEhcDVlEIQFpBcdHfWPujDXPw+X3DcnzLa9UjZa6ElNpqRGuSMRevFR8YMKtMWgXZN1L56
BvPjwY99FMxFg3O0NiCVKWfKl26XgfGsf5Y1EYtnzq/7Vvcrdb6IMJmHrUOsAebFKayaEkzTj8NL
Qj5+Zuw21dEp0grTZfuJgSaJhXPMjjKoOfvaH6LTdvHMt06jMiCaXmiA3kVQohe1gaNoAHUqfhj4
3LqgXMV8hNEr2/tsAm4y7tbbbxtTaGdAIoTBvYE1Lx/EQ9D078FYh0mQNAcTfCxfvWB/Dl3DzA8T
miQwlXnm06ZwYa9FyEH6oKQlDbWc132yfAvno8l+nglgbD/2OHpqigdHll+gxqftORzAcjcUXaXc
hp6dJz7k6tURX/PxzC/a8xqWjOVCaetBN/Vv8CjJ+OV5xckdTRdPEhiHrfJJFe1zyc2O7Detz7a/
xbi7F1lVtTw5yRmRjnukfWIBvylpDJu1kRbxRVU/1RzpSnokAFUe6BCtcS5aiVbcr8hybYa7+ORs
JRsRtgunibweHiAcK6nOPLOdVY2koCRsUMdLWE2MsUdM+ROUBOiYgjkqTLTMg0OSdKoeQwOm0RvO
Ih8gU9+RmgBS6W/YUZ7UuqRYrUOPxEzn4/4LCG8seSgzQVUG2+SP1rbM0K8L6jRNzyAiKcLL17cS
NoXZhHUhifJzO52gVG9nXRrCrbrqhGtizcYoehARigHWSeeGBN8GsbQS4zmziCurZ/akAph6xlfP
JoDjb135nhHbD2XnEeo0gruZlMxTzcdycZw8G0wYjPf2Z4qbONBTIBrSXU6ssmqO9ggRdt8dwAuj
6u1ZBs0P+6m9Vy7vdnwZbH90mjYkpJ7Hbipx/cgiXB6PCt2+naDRb1DvczWrSc/2jlqq/oE+GNtT
tcf4Vrvsdu+95EpDQH19KVzDOuKS2zQTj+MJLy5nC2IxKN8gQk60Kn6voaP2pyJXE9/QptJKe+Kv
te90cwizZuBd5F53z35WRoBHHv8bji3QAm/oz7g70Scrb5jMgalrBahXdE46nQ1yAwwrERF7yiTf
E+dt0JHUjMdW6he40HEfCF9JdVl/5+uD0HLvCGNQl0T6UNd09DWSaZ+DiT80JfI5kUEntpJEYoIo
3R5/hy+I6+kvimgYT0F1jiXQR2Z94anVmGDVjzu25P/8l//UK7Luv16dOCC4osBxotDROHdiZDLN
FNPr3UIsWsrnD+bi5BkvJIO5fSqE03MJfB5ablr24a4OMqCrEkruY9TgJLgyMRYhfbTy/EMadstP
n6fU+frycz1Uc2llWhQWFMAv7PmByRjDXpIccSKFejdx5CptbKC4PjQXV3BpoAq1//rsUqClMALd
2FWTu9y9u6PhCO5d2YPYTacAqDowO3jTNzJxtp85QI3ZnKFe/ZVDp0Rg+/IoKIqzSUIzvtSAA3zY
YDvObZyIzlS07PZR1U/7M1ZQf/L0JZVYnctXDsK+mC+em1WTF7T5R6KajI+jPf2hmrF/TgJ2/UNz
jOCNxCwMCCZwlDGzWOOTIRoKzOolbBjxHBWj2w9RODrGGF6nGHIGraip4/HBIIH6ZM5ZgQjxJ8jG
NlZnqAOvT9AoBBDVy3y2SEnxl/kjsHXGefFjyBrC5kHLo4PIvYGYd5c5JroXMOcOvNalsxdBG1w1
T62jKQTOq1lW2cmjJng/Cjt071a+8H/misDKAEQeNFlE1pk1QANrXDY6pbK5/jQam3ZpX8W4+2/K
qkI280X/OLBxkRMizZ/1G4StIwSwr6m8gNQsJUGeafhxJ2+ibLnUi9zaLyj2MWvwMihwUfNj0iUD
o5h3IQbYcTCkHHljCSVxuXeflFlEFwaRNBTnzJF3TrS3QzyKwUXB6M0kZ8fHeXNn9PzZtNV/RD1m
CXYZaTEJcH1Ee1Lp5GI5Eiu45u3cEayScZBtro2ZM+HpUjxejVquqD8tWcjf/TgdS0i7Lk2b65MD
Fs62EAl9ZekXphSvfvx6WsCtDMGj6SQPfph54YNpuZrLTPW8vPtMEj2oIIa5Jin7cZZZStNYVaJ5
PA1Ek1nwgSg0XRMtrmc2O0XoFge89SNLdeZSdNfFgkkhPcHzVkJqnDGVlOE+mYIdgu6GLB6TEeNo
7xj6B6Uew9/Hj7LUbeCTjnEkwTxsUnRK9eGTp2Y1CArRrMZRKA8jXLqFJ1sADWtjJIB6q1rVfFJu
iz4SjvSHasy8Q5TVAWt+Hz56XLHmd+WCK7xUqEpZltM2UoclcihHdrJd2JoLgfqMtUSBYhsjYOMA
yMm55zDbTAVqv6m7RqOhK5ymMazJw3hnJwjDhn8eoMehNbHnmTG0Ar/Jiq4905Pw8q4e6FI8DU6E
cdbKGl1xZ+JMfoElhZFkbSDCpRGhDS1DkOwGzg4s7HEA39fGRPszIcTbbfr9MO+pN2W8aFBoAay4
bhj7PYS2Ofwugu/sSsX23/rdMvIknzEZc8jl2gGh7y9JLB/1t3B9pqqo2ygBvFFCnwGbvsGgAmAs
JGoDvnwOtBc1fxcWhzVBmuTlEIDFddy6hmzXKqf4YE2AzsJbz6awnKBDmhO0t5Fx1oK8Vi6hebdD
GobCXMo7q6IY20HRXH1UVGMU0Qkz0usedkWZ5m/Wy92n1ztll6DvsLjXsb1C7PrmALIiLDTUCKXj
dclX/NkwbKz8/NaPtPNV8M4TBBsHrr6IpHcaukUGp1ThBVO2pT5yt0KiE/Ox7TacBC9UFstT4MMz
lYeSY0HT7eiaG4zRVLISiOc6ecoyJUIwwpaNO7gB2l4Kn/763eeV5uTG9UFyDl3jPVpKTZTdRKuF
LnJ6eazk9RiIa9S5KkXMLqbRgBrsOIpOWKM3sN92TtYsOdYLSCa4/PGnwnM2CzgZv0wTjikG5ADu
h+pE6wqSdALmPNftRmZt5WU8uOw5N/mKX1ix0uTQa4vJMstEQa/LX5dzrcXZZEruObIJH1t0UiW7
pCCdABpYELHtDNFiUnoQ0XVh1GUt/5zMn8QN8qjxsK3oqiQDjtrN8KI2vuzxcEtGXp7Z959oxZGk
AtDiKNBS9VcwVeuvOGOuAiWBv+EYy5OJRUh3UE54y/czfIQvl3sLO2FhojvX87iQQ3uFtWKfSuAM
Nfdv/u5htXQlXB5oJ2ybrJO4VEi30gLO8kMKvA/s7lJ2m5jwYYoOmD6Sy/Qgk1GHOBhY6r4m9WPB
j2OdxUUgod2V7Mw1Sem9qHdEJ9sowgFdqGEK4+aI/KjWz2SQJRLCchZyc79CoeR3kjN/aDO5wSPB
Hf4Gn1oBQ5yS4dc2xOjCqduFpKeRP+wGGexDUFKiUAKlAL9E0iueRsyIVs3ZAnZqp+jdEdKSuNle
wv9rO8Veydl+atfR5OzJHTYYy5YI7V09XNhVcaBbXutAt5bXl+vGkPfkm5IPwSLH3R3QIR1GkMNk
QjGesIP5v7zg0ZzPjZT3ZCNMfKBsrX9+Uh1dY4aMx26JRiL2Gq329PvSHQhf8nsMQP9lJ6dHPf6k
Ex7sZ2EtsDjSc/Vqqs2B+JmnL+iYDSgAjZ8N/KmCLE06zH74ZBFVQGQarSzu2SO2K2KyEkPFPYCM
9uEmIsVewpPY9WT56zRsSK8I22aPDj6Rv1y+iBv+s10beTTOyGX9w4OuP6/ug0fYkYDEffMugMAn
G9WEy77ktrNGVnptq4IgTkhjtZN4xQcRJEz7vv/udhpso7aNsj1D6m/Cp4uqOeKrnIHCs+AmGFrs
gaAmeWC25I2F8XJpqfRNW9c2oR37rzkyuMS/NKX4NeH2uDscy2zIUMcjypIkNa3fH3lMYgRHYkHX
ImCGoGc24rvTFSZ6bOHi8dnN+4KNhudOs/FTd9lhj3pJTpJbrfAz+CuwZRKhpjTHlwaAiDWybTBr
YtJOxyqat66KIYa23jZElEpMVcZ992bViYPbvgdszerrHaHARx5lDGjkGDDOcQE+VHitiBRMZMoR
nK5c8VjdaEY2ZLKHIsKM9p9kdISe6fMpswwWX1OyaRgRqgVHF9x6tjKIFsc8Kl0pQpLm1gtlHfxK
lhqQt8i/2nB0l/5Lg5oR+F5sNzhErFKeaw57M9Uue74fijFSfJMii8HoTrutsziQeLoJeyT1/qd2
TTUsZHK2eruTSJeawCqYPb+z0pil+8mLjCQR7M+tZ4loKLh8Egjuir1M0N1RvznLX4IAngyN5DEC
Efe53BA6gOT7qcenxIZrWVfsOv09zyf/xf92KpHdkdH9NuPeo0z3e//lLHVnC8Zk3sPzoKsmCbZT
dU61F1kNgcqMuOzRJGOIqOYjPcE+MSeapmsMfB6ybbRNYBr7kox30mPUd8g//3eYSla+Z+uI7TkM
RIVy6H+OIl2OqZltip6ndyoF+nOfxrGOo8qbkIuPh4JsoAdFADW1uLfXaSUfAX8JJY/ms1z+MxTm
YCFrKuhLsNxlzezWDE8poTvcPI7Q9QpyH/Mwl2MLauPVYLr8m+bHlNXL2Fww6V4+D4W2wxnV3zRc
2veirVMBZFMi8kqsMwOQn6UMlBB6CtDmML1Dx254Pgdic/R102hCOJCUJksB2+8JtijYCnkvMzJf
yLLOOIY8vevOKsea19yM0QvREq72xXhbV6o/saoPrBhAWHMPwyANUxl3a5jzwahFqqLDGLXGorWm
DJo+2fbCxeLbQ6gcJbrMzF9hFLL0LiCtZbfp9YfS7DveL12doS/xJZvsPI6aDfu4FjY6pPLJ1uaW
rAc+4rBm6RAJo607yCjTvhVMehuirTTayBGjSBL7so5rWAmpa2MTqmj0ZP9gkxvQvB6fL724v5hp
vQL84QakikJmeCZGIM88xmb/7+NPzEOeuY3iKwLuoXIISasiZ4gtNTmzeCro6gih+lHbjnYiJsDX
RzvgKIv41twxHMiJqwWaxkqHd6BhiQfw2jGSpCA0XQgHxto9KmR6nsr35QLF0Y1nulHRJKe4EgbH
NBr3pDu+/qB1RV1UUzenp2tRld8BbsZg0q3JUNj8K/iTSPFECFCicA6rYAo1iRuvnribAzdAZRba
Rj6hM5bkZh6PwNwLx5eKHvTbBWY9nR8RhO9l9UbMYOdfbSSSIiXZ5cD7Cw0+I6AwRqLO+G0ZtLL3
2l2BIhfyWp5a0X7RsHePflS+sPI4kDRQqYl65gKITz30u0375ZfHX9ZBc2EvFPQmUubD9Be/H9FE
v67q4mEmzfkamv7N64RFMkZl7h4+sYRxzqK9WwPiBxyR3wJCG/l3DsKgfQIbxx381G4CI+Yf50VZ
DrAPerayvB4xJsoXrp9P9VU5MheSqcZf0bRKOiryGPTA4BpkNnSLQmE5/RSCOie+zgvMPkOM5aIX
+UAyzgqQkksaXEoBup9CwjXpfXM+1RkhXJrxE+pXDjGLHJqAOYNltGeKu6DWkM9jh4ZQpaOrxG39
meRoWm8mhGc6Ow9dfMhV0yYWIzfwxFg3vVxspmlyUjowbeYMX/lYnWBhvQIHn+PEY4242qIDO/Xx
e7cmu1vYWnxjXdeAKoPdHI63iM084x8iUi0A9wM3Sscg7BEM5iHm5o5b70M014uS1Dh5EtZ42ly9
r47YBAchxUUjNZ6BKL0d6S751cao5zZt2cuoC7d++onGMB4VsnYxajWD89InVDJ0nYn6SR0u2cz+
YnM4TIcJY8xejoKY8IchBQI7ao8gii4D4G67mD+R87wT7f+3zQJjDVnf3JMggnlSMCGpoPXostmY
5fB8LF3svNBKMxJBlsvqLyJo+Lte6QxxxeBfFRwlW3a3ILpnyDC6LNmt4T2davacnXRAvx1vl/Rw
a9X/sb4xHiS6B+wnFhHeUDiH6dHaSm+4D+XrBSawBbaaR4cCCPEI2RMVus4QCyfMzn2Ki0mCuBlf
X7W7hP54TN65/hf6EcDjc0xSxeslrvEGiMUzmm7EAiISrOB/xHGoiyxw1fH8+zNkuDkRaAFzeE7X
Q1Zdrmb7Yb57G2CurtHjbpa6Pr+jifZmlSJggvvxg/kBJVgOuo5sQoEMnNAdUOd4+nPjskH4xV6R
wZEMEQ5ezH9Yu5ezb/YOgONXkK9BnAG1MYfUq3u4Mf20ofsmQMzPEl/BzZdlyvWvBakMkXAUvJfN
uFda1yYV95kIY9P8u7TegdjIEHHtjZXjttHKyctjeujh1hMPgfVtREkHT+sogNrS7sylX6dqoaAM
sWAPHv2Tf18UYg5NL6VfQBxnJdWXixuQACeX4TEMjsvgggCrbfyQzYLid1AiILgR8OP9cII2Ea1E
eJE7NZ/uZz8vCkcjhc4mEtZtlRAnygKx/OwRp3hl3zjhKWvf/CroRecpjgiI17P2dq+MuM6WRwCT
x/fpzYATIEd4BXI0Z8oT+UEpmB+xyq8R4xYiwCka1tJNKq8qrMT/jnZV4Ns3/vkjjMXbA06VzAld
hzns2UyKDTu7Oogiu9Ukm0HvduniTAyeGqKED2IeheUChWs5M//P39C3eFZQ5LRMu27s1ZJnOVQg
PQhDrQ8ZzIkg2ZpJsSt+Q0oh/3l8eYfBzGlB8nFZAcuuCk9tVRiDD5yFkUvc/WgVdxmbJ31liibz
hpEacM4mmkJJdd59kqB1d45xhsJghgdR4mkOv+Z6gu7NNmyUfWBnUmZ1eDE4wkCLnGRVyuVVEViJ
V55JK++e6KS4o6IgxVbBKjV0ZSm9mksM4q6hnKQs7/1YqckGo8DuOIfwhkb7rzXTPvZzbdgwUQz6
BNrNQ5gqhxGRc9sVw8hJ1BXZlLYvOCqArNOScDKFBd/JLolD/SX9IwuFi4EXey3sa6h1Ay7uRcI8
C7qj/KXHIszq8Jjrumx0LqmOwsFfAF3ePE/KttHYZ41aXzFuGUZfLQ53tm0qxoIUYqoLf46QKaUM
Wp+u/MewKsGMEi1FznjX0hPzAjgniJW4Vq9hs2oRy4Sm9DETpIgEZL7uLoba908dYGRfLBOKymxW
KTfrpmd0xNcNYp4CCk/LjbiXQNjvkbOCKiT3Dkzj2zTHozUdqh3sSMvLLhT1k3SgJXB8LLPQ/naI
2uhmxk18lo+IHmMnxA1GpaZEeblGbKn86jBLflib8D/PuFSof7eAoUfXOxpX0tweOQ3mTvijoEem
Ee1hwdTtLVLyNsbzWL9l+6OaBwuM2svKEV3C7moI7zGeS8bOS4yLx4BqrDLpBpJ07R3nDPKxTLyO
klwq6n25/w+jyM5bQFF2w/HWRyVFadKeECmCwV33FNWBpH4mSEdxo4l80BuBZTqASk5OlhyLWhyN
buggMHjsGKf4mR24aO6ySi5eKlONyQKssM7bz679XBNLW4lAxQWiGZNXKxS5tanptK0oXUKP+scI
ygt5cMlvfFna4LoKqBjDygC1ZPDnnhkJv5HtU8mYOo2HVg1Fzf17PiYHZFc053z+zFkt1LgKtB0J
jgQvDN9R8o+YBV3tFGylqoOD2ZtC4TsEU6EZsj5pn7c+SMp7FB3/b3LyhdeRcM2zolTNVIGb2VIM
1JkAAcjU5uos8o0wqV3aui9Aciv3fhv6SvqmdQyE8l0UdPyeQgTYIFXnVsRJJzhsrGqH0GqehnhS
AIUeZ/YLGGOuRoSCZGdGH4nTtIPYy9vPkhnxQ3u9PucaFYnTrowD+5yCqcBFcZhRiL3wMoG9vH0n
UpFtnNx9Cu5HIfe/GIFvTC7rzD5007xS+stvYrwWJnnmNiEiamX8f2wI1VVwEnNasvg4J8Fj5ThH
7sUhXylDXpMEOB6swaCYlWsbS+jIOb+hs6cTtyS0PRWxEwK/r7xWVwxFog6CFfJG+f8BXzL3ipxe
dDI4nonYP0atfSc8c+DVmKZR6FM1Ry8vJIOda/37MOImtGZJp95ByqtYJkY7vHrl/M31SOGTSjrd
ow0cO3kL6JKPF3C3ulxUpD+UD2N25lKxBAVibk0ZfIV26cAChRfqrb6JPwHnQ/U+1vw7nAg7+mY/
1d1euHyUp6Iu/1Y+g8AEj5DQLDMG2aJ/Qzzuo9u1dOFgdTElNBkvOScB/gKWeekpz8n11kGgKkPt
bf+eHblmQ6Z0XSSBZucsouqck2SMjnb6yhU4wt5LEtJ93J+FI6pOeHliSiJvZuk7LTt9PVdRxw9D
VvkVpMmOPk7QItPSKdKM8aMdFBUEDR2QK16PIxZzGO5Ls8xPMRo6xYG/6NZZ08evjo5rdgdtCBY+
7fHhQlqWBE9acfEMJl7kpRdNWAS9AUnvQOm8ZeG1jsPWmqbf20qfmgGQdLUFO3oph4/zKAQZkzam
qpyZGxvtLduRhZAplEsLxGLAexu9aGopAx//CihByIta9D6b7hq+y00llB8T3rH1Dy2zmnsx+YiK
XEZ9qcwdLpw4WJjEo2IpOaUoPuP5bTMCjrkyZ3hAvKaqWZz4AatuzASJnP6f15Lnii2liEilUy36
5is9gph8UHI1oUpt3YKHufaV9t5FnVEooyGv5eXTGcpGgoV/2WEqGHSPFK5qVHwyiU3LW8EZiI/M
32ObINkoXUiH2Gj0fqhoxqQG5vAiVKjIij/Sw8ujWf/1MurDemWTY+lO0MUtjBR0Lwezd/CPAkkK
j5xX7+QqGNMeSPfeodY6PORqTp1A5+SAaLziyz7VtnaXqSOBK0BLa8IVMHeo9eIPIiSPkKQHEfO4
Nbmq6yuXQGiCi7AOXhqnHU+/Fv22Yzz9gf6m7c1G9YPK97pd3PccNIHarr7gZAOUG4GOviEoyamS
gSfS2Nb5StQ+XAcIyjvAjX9GwaFT9JWjduz4hO3PlXPfphFCsea7dJxWA0UuzSAusDWKt+l/rJYe
N+aEDqp66G6oqVNsQqK3H2jQOS7kb7aHoIVsEX77Lp7K+Q9xtBfegVsLLi1aW72P64f5RbLs/LLo
6BwLJOmDUjYy+yP336RQclckBvMgO7vf+LEiB+hoKTFXbMHdR1Z6gkrZ09vLH2u7nAPNBzIG9sBC
B5WfcZN7mA4ZvPt1SgSZsQhVJvFFz6gAOf/ePfGeHHdE210XHPHqUDdn03/j5TeWsg52exJLU6kJ
k+xC2BWvpthy0GlBUqp7/u8h+l4SQ302GfRoTzpFVToYR/SLQ+qOSgz6A1eFaR3j2XPUmpicYshm
8khkWThDlm1WMFIFDo6oGeT+x//461yoesw1UDbs9ko61q52eyqnKXbNCqn7k6eYXNBFseO/7W27
p/co+G3LfyOLoPU5OddHJ4rH+NnSBG0pd6hxjSxLAXFBWWgnyvCh6onTiNDA/grqjUlXDaJyF6kh
V/z1wmCHsTo/ioQ57OOKzNMeJ2Iy1ROkup4uLn+RbtWpVFH/xD735ctUYSHAsrmA51gMDx8t7goo
GZalIYFFGOT2GGO/BceJhVXiZUCa2ak42F7srOyo7y7TlHzsB0YThaW6v8V7aeMBQdoKeqr9bxpb
Jfpe+ZbDM8YxxgUZ4L0qfhHf/eyjd/tt5gfWEzRwfv2cHHZaozrEuyLKJ/u/9j1JhItYx75ScgjA
7ghcVIp/2PE42IKEwj3kukm47cDHX444Gra/2bz12HzQrU6Mydisc2EUcLxVGSB51WmiX+JuTXJA
mfChZMipyAzLliVr6TcjdHmA/BO/KPrIpBSqFLoWqFHXhH2yWETrvlpSzvbTqdMEcv+YFkVJg7su
oQ+cRkw3c6nfJHh7whizfFdpQ1FApFts0vVEUjp5o4rwnb5SkELTR7POckcyzE6hLH1TrTVrUvJ2
4jQ7HSsRshxDWWaLOZX5LPdgmGY4fUPMuFXLWvJN2gZrqGZgEcLQgwd+l3NBA1CcDI5fyrJ3V9fC
jM3kSfEFSqvVYbROL9rHwYKrIUR2HsBX915csDUv1E05SANPWKtR1yFkfGv0/O2ELt3Sp9bpENak
AXZ8v2mntk9P7AluazbynL/d07TNZJNdqeSJvJsCgKBvQPgdLDox3+LAHxBkwPCSyt6mRTMqUayF
nTV1MuZPe0URkkMyjOY2rtvIhmY8gnl+KnBQ8A4tencpllM3xNhYKkKWFZ02m7Ge66bwEkEjMbv8
pnwnD7Tm0tXqP+QX2IsSpGH+n/41ZHBe7FcDVeRV2s9HMia7++L9XlU7NhKJhk+Hfaxe9hpeUIyE
QJ7ohNtfBggdoU3U7ltxLdFM6713jt0aa17hZDojsY327OvF3GFvizghRQ1TZf3AkgcEPlxhssYS
hs2YfpNPUaDCE9Hrl1Ki37e1d+xarjVu1N9RvCe2GykkOWypktSnhCznjJz3lOV3ad8AYdA6CEgk
zniczP+67wS2HfrQJIhv98W7aqiXvPHDRTEW9pK089/Mba+1Ntee1b0T3tcbypU5oT+gDYYvMftZ
HSoh8Z2aAehrQcZyQAx7fOTV0V2fMBpDDyCiVOcj6kvtR/BfnfdVJb13faP+YATLkoQQBvP9lIJe
XPmtrnc67b651zB/2cYmu7/rv4OpCS+YPJH5EYuXae7UnotX6tvyowsfl6HJAAqVdhK6TMeYvIxb
yng0b0fl5lSVSVPaJoKHSkG2rvLFtdCcITEKsh/D80oJtJihNpcL++8x+Ih2qDVx6t9/5sk6lUbj
XP/e4rDIoUnhSSPxLJCZaA6aWfc2PV52dzzOCbUcYhnW5gqdsMcN1M265GpXR6ZY7CSWIyAwsXFB
JEk/mmCPiuQ/1KKz6fRIh4XDxLSnwkF1tJFoXIYFO/qyA9ypGC/orZ2yim+Jyc56808E8CtQ3f1R
WY7/eBln798ZXHld9fZ0q9Olz87yqrkz737T8+FzdVCwf5G7/dQ6HZx25uyBbt5vTX7w7J1L1OtR
SdlbqsdbJbqGVqoshzcS0JD9G8Z57RH5RVqh++2Qjo5UFLncdXtPTKhdMIDyaWasT8yHA/tujpT1
Zi1mn0LWcfXjp/rU0COZPkbmzeDpiMx8Q4yKE6TcIFeaQ26iDbWNSu5hrcPLhxv4JMfJOVLgMrLs
aiKygyqyIEP9A8m5hTLAcQXDHM7ilCdjQffwb71XoPUWbfjaavsLzomJgNtWis4KCi551lANpu94
f8pTr0C/xsQz1BKTSgq0QlXLGKrDubS1Uf8+Y4gMLdsw9Bfn7+8bsBeK9el/Ax8easNI8QVtB05q
3nycfCyrQjDgEUAESdwM2AWuGAdg9oQ8svKWLwG4+P1Xo2jL9YuQSxv0CLLIBsOIeAlawrZ6Ltgp
25ok7aNF9MFA8Yq3QaQDjvLBgVc+9Fh/12/cTrinnFdQ5/pGwrxjMwODLj9cOG2YMGq0HBNaUy+h
6DBFDsR0heLJ94uK613Ha0CCEm68jq/8QiUhJuWD9pVWoTxda7NxVNlfK2NhCQoy/z8oHWvjHZKp
I1qYbOqCXMWtQNDgRUbhUKZIYUa7RKTYAdUMrbS6Q+L/dAUSKDBspXNBwNVnMrqyZer5N22fnZwm
B0SRne3YU8S7zlG4mHGynLreMgnLmLPb+Z8gAGnYqEh5vMuzCbYjf5pcnU+xbzVpwXf+0VxFY/qB
yO2sFbub+lf4CXtKvZJoB7bH7Q3QfU6Fnkm1w6O8XdFF0BFkGmlTSVa1UyJsTxKktSO0KxzmVEWv
8O/xTdhtDBp4v1VcU0c4d8eAsscTafqWahs9P9kG7r+07RQA34v/rz8ehXo9mV6i0rp+14NjZETL
V4lpXnftG79t89gSmK6JYB4M8agc1tL6j8I+W9za8CwhDR7vTKdxnFOzBG/L7jCm1XaMIKxvINk1
HRTJnH+JbKLchbcou1bc1jecLVFucbKXLZyN3v1UkVfyANuflGLbpveL7KBijF+puh4reycVaZu1
KGcuJc5nqBs5Jx39FSFa/TRQ5LqnT5kOKa58i8iMunQWsMtHV4CV3JdmUxUDMy9/2Dmx4HpD84i5
YenKH4Mz5pFsmEA7Po9srur2giRusMKipd6nIUssUulpAZK/xGRgVpWlVwzawt2UAkX+hTxCA3XH
w6ewoeqxLn/WyoOKPSsyR8mEiCMk7PnvldewJauWbL7BDEELGpzQJaoM5ShlxiSYGkRfDlaukL5f
evY/Ts0+FxqzruIStupwdie4aFZtHPiyND14LH3LVLiMo9Upsi+geujbmbC+i0tWSrilRYwkBJXc
oNDxsA8yvu+6xAr+4iEouGw+AxWP/2aYx+J8UCEa8MHpBK08iKBnRRz/Nc9NI3FRX3BTMpmGJ2uC
dA/UkqbtgT5UYs7gMAT8uenF2VKtUepV5ZwsVgIHda6Sbim97BgYZHbkVvl+amkz958CFhTsy5ZI
LnTmbjWdFKYh5/1LuC5ebbSkOZR20vQuZZEYUWzIc5on73uGiVdbMSP83bV0akBnuWs6jZz1yXn8
VlvPYAvfFQXFoJ/m3v8uv2sQRb3d8f+LwxCFHM0A4hpbup9ZHfziWFpQB5r1KAbiXIXzWs5idQwg
lcsqroQCVF/CGeZxKX1KZtF/Rge7vepLWoDkb+Qm9AxuVND4+YLZZy+utqJN8on8vnVFJyY/cE9a
UGOy2YgpkVGT6OKYDtRowzGOjY3bTvO/Zv/S6mBLwYM5qKKkgrUs/3Kt7aVdYB2UuilDqqNjA93a
1zypswgRLwIOiu2s5btLZUlEWq2RtDoljfdEdceHGvXvC2XSH7zzkw6si1JgGj4TaWOhyE+xF+VW
i+IOJ7dJxeUk58/phKjaxDETgWnbT8Gm+/vg1JzkTS/YJJsGOxpoJakTeKyABbFjnxUTyaFYj80W
78nv4ycP0p85Z0F8oNbIQVRbjT9osowxKWiLxv7ZlHJK2czyc92cNmfBDkOi00kMVbTT/aTa8Xhu
u+BN0ujpj4PTXP/U1YoZwqfbjpH9s5XdEn4HAcfdRFyu4P3ld2P9W61FDoEhVmYRxtZO/HVL19pw
/BJvXAlko5XJKQCneKYb5fETAXpG/6dz9m0H80SXQjabRcN7Hq1hVyuuPLYPaIp7lEpqv7ya9Qap
hHE+e9Yf35tFKa5P7+ZcOtYbMJImgifAw3p2+5dFmC1KYyso7/vXWRH/obdTU0Lu6HBnYz05ws5z
Klj5KSgqql9BY3HilVj60Yo/fGB5LWl1YjMZ+Jclexm52Y/1DYIuJam8wVLpqgyaVCPwNtz7E9OV
MaBEOM12SqGBnRk7useWKPOi2QfKjb1afhbQDWc70fmvWPOCvOaycQHPMtncV+aL8Yuzkk3qiCql
Y92d0x5NEixa0azjREXzU3hQF5kHu6LCzDnHnVS45seO5RDpHPvRWJsNGnx7Ha1wEc4HpIWmzMDz
c2Dd9PrG8AgiljPErTwRXVlTERhE9yeas1mSLQofmz7JX90n6Ftg51IiX3Gp698hI69is6qdPUNw
EU44keOsXIMY3ZX9d15bRlsA6eLzr8LrbP7E15hL5wpTOHTNZOOY2hdCX4buVS3LcG5f4rWIa+A/
8t3Y/jPjAB3DA6fIQImsjcXS2hqVsvr0OReR/jOiY19viUzQU8jpu/H1dBCbL+jTJLEXx26oQRI+
wYlivq4qHoUNztCZ8hEq0TBu+C33/NeA5xBKX3ADWkwgjjlYCaY8ok+uM0AUQGSNsRU/XBSZ8VlA
TS6nc0vrWjMj2NhnKq4JDXIl5M/76ia0dzGgsUHjdoSjBspm1PYdfbYC+JrzqJxSNphYhldQKhrp
DPnbEMLRLJ967jgk7l7I/1mtwY3OT+JNjyO9hJwDIVB77YY3uh2qlrlMzVUYJ0m8T/ht20jD6hwz
NVmn3IzPfACM6kI24EfgghxW3E0HkEtTNLn+cC6MBVY27/jrIT3YtYNwdZKVH0k/Y0Js6Ux+A1p8
ZDFwH7PJpO9Se8C+V5UbAIEPi6nGygGR1/UqyY/xrqYeTzcpBbK4IkbySev32Ra7mI5HSRc4CUo2
2wPZB0QJSPaDf3cVrYhdXFXP/tDTGbbFKyB8LovejYvwJWDExe/fgoGwRR+fFXm7f5ELVkVxfP2g
z/5m3jr9eCyFLUL4zXeaCfZDri9KhBm2p1MYVx/UYdMOgnNbu3UnieriMsSuKovxOiXY2aSS8MHG
7/u8hOJk5Cf3vP9tlDakHJ8x7KCk19YUxMgPJ+nFiyjz59skJsmk4fRRY+bBAizZS3PsUAgrkHkS
dfAOFQGBF5ivUUEhvY84SbxNpRL4RJB8UKqy4nZYOO4dTTXVecC6tAszqzmNmTTiV0YPQQF42PXG
NMsLy8wfoFhyueTnDY2ZGSS2r4q946MnHVM3fuXqvoAZ6EtGbKtsvQIj99d4uI64Lg/lWyqaNrOz
tDotkpIj7+3vwjb3PcYvchzJaCx7bX6iWs79+fPsYNetJaDYUW95Iuo0TsprB4aDsWd6/pdPtqb5
XicMr3QdQH+qsm3ZsNFjIV9RjFLK/kIgKpfsud7MA00S6hdVjCyoutw2xV04DpKGzmNXMk63GPrU
I8FAbLn+r2CHweq4yfhvfh9GqRUOg89Nh46UjqTFidvNe+7wPhq6EbbxEgm+oq28KoUqY6IVjj4I
xZGEVXjs3jQuVlahY8LKBC2swTLtiFftVIDNLDevrmKt3XKeTb03G7lIlvzGVapOSvVllDsUyTSn
zrgDwBZVMwulZ+mrqL87KI/rha+oy1TNabILh/ukOKvhseQb9387lxV7z8effpIP6CouhnBMfcHT
jsRhv/gYGFPJ+tysMgYXNd3+b4p8o5B7aGvgUWZpdSkDzYc0qAlciWegqDThSNQMAWwq3HkKugFU
CpIDkkhA/HvCKiJER3RBgWIGCyxOJDcLMdzW3p7I13w4JkcIKGwelR9XPJHJfe5nJ7NrgZ77/b2M
awOAULo0zN3qc2V2PaLHCpR+nepVWdHUJ6ij+P7dBwU2pwASWBuWHiWi50L+tEOWJcVc0LLjImjE
+p3+Cbs0p87yKI59yk+/9g/LfprIKg6SkO/3QpxjrCVell4icq3ZP55Wx57K+NTPD41xHQnzXBH8
YHW5L9c8K5TMb9bp2wNTpJFbWvOE7WMkPvMRVzDFVB5d1AB6KzRhLtiPLSDEfxkjXknerZcEaSdG
sillWge9o0ExVs/qw0htgkiyGSnewE5YVryYCURV0olcpUCEEn/RQzw12wUkedsBdlr3MUtUdCXt
7tMKR8ZD063x4REwtbS1LtYqpktydHCE7cCtzIkbEMEiOIOHr/HDecV+oa2wfY/Hjd65jSSXmAIB
4mthd2d7PC3fiXjz9gh1VZ605fHtSCacdyncmU6fBiclFQagiRyhuwq13F7S3POIqpsN5qx2P5Cg
4YJGzWfZbkbI5pL2IUBNy/2XCTcLh0Q3Mk+KAeK5aJmTQKeEJISaY4/mw1KLpyoB0BMXUqVf5gnA
owyI5pxN8qC8LexnkKE65pXsBqRZZpXg+Ig2ku3uGtJYaC3ZCqTH5IGjPYGvsZsjQAawLB690LDN
Fy/uZSrblGjT9KLXgh2N3zOrXtHzdjhqBcXwQcs8FkmPGIosm4ZYtH+EbcSjoe8xOgwlg7NxJxdm
F8cWAgLb1HaIfigiAyn6vHpyXkHAW8o7fwAV2XWC9YqfRxkdgBW5C8V905NIZPiUCjGAEZARSiMV
Yk+XM5kZOXXr6zr6IllsvlQkC/P6A4bYNAg4ukSUCOrb9Iw0xOWByi9I4WmonQGoiM2sCHkAkJRg
ZbaZwRD70Ar40PAPdQr0HMoKaOH0rYd1n5HyETI6FPgVpBik9HC9735lkVdlQmsHHx8vPLLu1EXZ
br6lHm/Gmsu72er/9HWaTUmtA8E8ySsKHCcOd7B4EIiBhgXftkF8Jc5DJxQ1Rl+w/CszJ4T0gOYP
nyphPe2XUM7pDo7L0q75JpdQUo1bq0wA618Wukko6kTetkg+Sul56HQK7OcpHp+UC2SJzsgIIQBb
fUqYl/FxUQ+8SxPUw4lzUxrB0F86cdgMgGDDrujReOpDMCeUy0VeQfVl0q1OcuAbOKqvFzhyQREf
pqQGSBwVCBcOaiERyN87qzIbSZuJKy4NybHcSAMW8rl+Hze3HPIcRsMYRuFRpEXEwMHPF5LcYZqd
MLx8mMou/b3pofCc/P94Gf5gsVN1wF7/ABl7V9nyloLb7yjFjPWSZAQVNF6aeEjbvvjoaWPezNFo
3t7WTGtTTpPgfcfmPan1ebZve5WMaEi9o9o60Pg+DEtMmwLXBlYQ4L7kJW5rPaih86bKZIy2iqT9
p6aOiKnczwCWmdX87Q6duS7OYxQIWcmsXSVqythO1eLLtawNi8ClnnJsaPbMCwCIyoyp81AFGsW4
n+ErY2BwsfLhXjPf7K2LD1nyHfWSbLMSli4tJ7jHNQALu71dzap35+MElBUjcl24uP/34INMwO0X
SaU1dXRuuAvtfcnEhqaJ49D8bu0TLzqZihN+KxA5EGNjAJ4zYlXuzjDhOzUP5BVUp2zcaZZcsLMN
MzRokjX4CIKJIi6n8RQJzS43jUn48TLF9JCRwmwmMeFt7QJpvvOp6cOzN2Z93nYFJl/lAmKxTKc8
YeY3ngcCI9SDWPwUJI32n052ujOn4nrXGfjlLFZQH2rfIkRYrv5LddZ3bkIoc8sJBXCb4ur/N2z9
vURlJeb8o+/oyg41PfvN9gAiBtNgOxK8M21bN2WQOjEyCq/ySIdEEnb1C88trB1StleIhXQ51MBt
d2j+G6Mp/3HhB2qw40PMA01v7JmVyEnYYxM0i+w2gpsPBBsbQ26ERUtJPF93kSItCOF3J3olS1N5
mCX92WcroUiMCOwiqNnrzs2z24WriJToFCcR8kyVWy7U6NU+Hqi56P2pYHKVBCEpnHlY+bzTAaTy
ufsHAes1or3m7WR6NM8NVvNulx/2pFknBdwUYsF/uFK92Fkn1cjpxSKPqb2EY9w/rUjjdVRQh6ep
fWnG2ggmD433seoTjLoZn/v3dsUPpEmrs9ARECbPwbcGesxpBV+rojq8EcNaD3JhHFqFUJDW4u2/
BOZ3WbRnLzwMclTx8ARhPjVb1FDxEKHWp2yAdHWBbv8llM3YC3aq0wpYdPZkG4CbjX2mRokbn8qR
BBPFnUgJlJXz8iGX8zSYjE7/+BK2IhWlJHT30lOdLHHGQtx1jS9llUFGFxAqr2gi85VRVxJ/kBh1
XCxj7gGXYq0+uwJ+WX2k8Y+ZT5GJQXLPQPGvaGceGPMMWKcwAEcRQl9ep39zI+Ehiwln2ehbwF+5
Z0U3hzZL6/95deLoSyZ3B0ZCEI7Lx/+o7OL9hEJOVaEI7aaJAltqh0438vkKL6jQcP+bFu9GkZ2E
t6cnk24FAe1ZmR99GwR1yEote+Z93E2B86FJQY9XAKAAtB7jvMb/9/md7Uhy//eyOVtEYrYyuEr8
/q7E2uFeqhn2rWLQLxQLERhMSIfaJRi72lmvdnPS2crLUViZbe9EmmL373FfogglMARsr3mXaBHa
dV2aFuF9S4e7LHI75KT8F0KyicqeUBBu1M0PgqUM+PXdtfjn/hc5iF/4y9zUgQQRdxTPmk8q2pRc
YYFv3DFZRtGDJx1qCL/n9yk4jTpOh5y3ucLNg9maIdNAVSSLL2VUibegtzW89wShSmu4zb5wIzr3
jwCc9gYHhND7aOOq06kqN89ihoTri/Q8MoCHr2yU8NV2BkWQpLlcroonEW86Hw/4/iZZrpZm/Ja3
vlgSy/wxoIrOTyoSKoIzL6QuJVzlDaD7/Mz04f64uAKPct+ZBDiR62vi2OQVm7bVsErEhJ1hafQV
/XfuQ0V4poKKRT0DrnOXZvOuVBwZ9OSIOMjv5QDTW8HEWPSywBw59U5ecwBWuXD6/AvuckVNDIaD
a8oq7qO5byJb7RyJecr1LPJ48njfGFMQ94A28SSxFVqtk0EJrjdd6OWPYtIwkxKRp+2MP9bjHC/d
V4TNm9stOSy4vS+meGGHCpZ9B+i0ztlTFlxtmevwExpsd9FCXBDqjZbRK5QA8RQwnagg3hbK0lcn
MgmDXevfrLruzLcrXSurRsU+NPZlen280eDLorr+tKt2mEnzu/DGp2G6o/ZWa8pkQKo3NYfGJUEN
Iw4GAs4TPPbM9bn6lho2QPFhV57CKiTkrKNCyD2gSMG8XnxkaOYJ+R1dFexNnF0limmkonbrANu2
NDYoJ0WqhEJst/7ciNKMoihTeddI7LNshiSXBPDTH1zKPFGtEfrSLpdIPhvRNzIoNmjnCMJE8Gb6
pHRNOCAExugY/xXzy9IoU+11piKc5hmaODF3iPlsMtw148k3tTtChrTd1rrTRqGbJEuD/MfdZFHX
CZuydFh3MVsBw/YCOGc91vKo21/NnXvb0itxvQELO4m9gWRhJfUc1WJmpL0pz1n2EDwRKC8/IIJg
UV+sM9+6aSGwqdLeGlSLnDoa4BwOXVnytN77NEjVwXG8reLrKZIGoF6ybUEawDJcrqn/XONum+pt
FAnvP7NSDSZu01ORVDF3MpAu0NJmBWWCBAZqmRuJo+tx09kI3y9ooR/RBRn9WYnMfK0LvHnnsjrY
8zPVQ75C8d9hxGeAUEDb7IYsYe8ptyQBn7O3pdt4I9UiaTIVNHg9xo9botk8qQcW5vaNYTWTx8Xi
DZvFncENPm6QSF314nUMirsfkJsofiB8zqFzNgwpH8CJGUoDqxyTm7YoBWh6IY7nfZ6wMIyyHhFu
LLkDmH7F+bqH2MzEs/E/7oV3BLvHy7sXw8gSLQ8B3y4aWMU24Nt3kmyN+BfLz00RyX+7288o7VK4
PSGqscSoaoaErJMwfxZT37A8XPJFOzZ6ROtccBlxrUm7naqGPhuM9GO19M8yQbn4OCXhqyYJolq2
BIAYSiONw2ragVUKyg2neMxAbnYUuCaTHjX6OHNtK6UDHeQyjnaREY3YykrL/Pklb5Tcdscu93Qw
mjUorSc4TH0OWyM284rrgLHjdKmTyxC0aMAJp1CVn/kvflKweWkRTZQhbo6cjBrg/TnxeHCBxnlO
reEVyfWCp5APZZPIBDY7n4yHlA7Amt8zSw/fF8XqXB7ikU+oG2bkeNwMCGYaZmk59jM19MBvNSyJ
ufI2j3QkN212ox4p4K6P2i0mLEXXVQatwMqzJ9L0Smum+2BrpQes53DT2woh8GRq5KnQut039L6b
5ROpGNUSjqRwva1H60nBTiXffWiJhwT8WX5bNc8VOTxMBvuEzuZZFJ7XAsfsfjuJ59A2IrIP18U9
hFIFHTVt15cgVk7RYYiLt7b+IsRo/ofbGX3D2RFkcd/9DLZ8HADWtqjT7ohk/kqBm4TksxRWS92R
l6oN3u9WGXgRA03yUrTGsCx9wD1tT4/fw69FF5zGwnce3TuZCTV2L8FRCLo1jh3NXswCmT/dxY2T
kfQNSsxSRoNd9BBuyVXh+51XAsWXwO/wkaIQVsO/Q3Lx61oV8Rh96/tyNUXfx5/1NWM1fxw+9WWJ
nBRy4sszHPuFBSuV/vipNn3X8UaelJ17b2AEc6IyNRdtDHuxSqG+Dj4JwyDGNDI/tIBfYeB3hTOO
6oBNEze0v/6hJ+XbhWq6DfWnEXmExS8Eqjzi56p2m3QKTcy7KAn3GMkVEV1fKWI/tmfM5oTwRGvf
7PEV1/VpzWJnzmXa300qgv2aRJP+FqbP6AlCYcw/B7jKogXaJH0AoKoS1Bmht5J+Y9id/PDPW3Ca
UzTp3CZ8kmG2GNVUne5JXouUejKTQiCn/beKtFZhM3WoMMG+E+lwYA21oiav4MwqxSwY/dHYAng8
hBGtvsSZyGT83la/y4vYQPDYROl0AOIJeU0pVkxLTP44ZWcjIoYRZAg+61++v64gzb1NNlnfc5qN
MxG9/EjrYftzlCefQYbjKdItl77kc0YydikuHFljos2BsElM7Yt5PlNVxV+mxD2xXNdQgD3AGv/0
0TlHal9CQwqrRP3KGkwxDvfNlJkRa7950k9D9rcnE3NLunSWQAMszHsxXuZDYTDULhTfQe0eU7s/
SYKBcMh1XNEnq2OTFIj+R3sc+OXnTfjjlE7fAgoqu7pR9A1Y8yKsauac0m6K4ZdSbscCOGXHPIl5
qbllUkwYF6hQfEaMJS2lMl4e62lbDbhQYLstDc9TDAu3suxRpMidQ/b1F6y+577sNBPuyTXq+et9
4FtG8BrKuAbrdq49xIhi9kBOg24IrAgkPhkuKPt1YlIQzQR598Ef8xUrG/wYXFB23wbObMzAm5I1
7yFzo6wLammz3ZVwva6FkG8M3Ksl3oxuofdgtKyu6QnVjJpcD7sT57RIF8yvX8KNLasW+oX+rwrE
aeOe3zdB4oE7zBh+t+Fd0Wg1lxhdPI100GdjJfoJOwoPxh1v8ha2w6AqJmfEizF3Ekz9XhFwkh4m
GV71SC97oNwRfU5g3I55lpbQArXeCTsQfK1jwMpVyA96kre7EEWnRF64CakHOVi9/4kz1m2gOxS9
+wizMKMmYMAocSHw0jChNlcZjS24O0Emh6TJRqoOwtRWw4r0wHoLkTa5ndGZk9QCMkxeUDsRT/uP
zcr1jtj3EEz0kzKr5izj6zqAVRsMfBzKD2ZiKOtr4Q8Pr9ZnApo3+X0l2jqvR7WeVKagvEDVfrFN
8AOeYNx/oKjQXVvq9DpoAQvjW9UUNEeZtCrVzh7gAmyNRJzgaV8BvKmw913NOAEUZNdfHrRpEFXE
sZUsM/lObTlqoZmvKgL0EWHvay3XG+s+S8h6YiyTl9jopoe3/44OjjxHY/pFoC7yVIri0exJxiUG
dKsZdVan8w57NtnwI6+O3e3vy//ABqk7zRiA+Sq1Az7vG5fCMwhVzGyOa74up6+wZa+RHgma1aX/
WY7URrFjtJw4QsyC6VpgM5TcimhXOXVO0etsAtVVOHyg+Vn0unA1fyka7mlBDcwrGuj6zq/qYY9u
NeK8GNghbZbgc6w/PHdvy9Jama8B/bFjKG9kGsOv1A6imsQoOMals32ZdJRZdFKWRQgXLqYWc+ZL
HX5l3rMlFTYtKjp7hR2a6i2M+nhvHvB2mO/3IfsBwQgU6jb782Dr4V3yWGPieXri295l3GAvdwRD
UUGb++feP0xwHGj6RwXgeJ7tyaePleGlSE/wr9E2zGri+Q/5S904BORXO+fDxQWMHFxlwIIDOAkh
RH8rIujJyFkWafRYrt0MUtvCrxA8LXTD+GjK1jE5pxeEEGjejV3WqDGq49LSYJEOHSFLQHTz88Qc
s98UlPnVxQepzb3u2mBkNPyay8RztxwRQXpc1lbge0Ukz2DLmhxy70QTivJx0VdkLoPuNRt7KnG4
ZjFys2FwzhygeL1lgCRoeD57WgNcB+CgGBvbF5a8ege7NU6rrvPxnVW8pkeGQ/DQPnmaHj338nWe
BYXkHudqVslNKp/xuyNU2izW/UM3+iqanzkARzuF2Jcyr/6TtnPf4KNLupvUUDYdzNoYT8cLi5H/
YAOUg9OR7Ogj/wSm5M4MVB2ti8k52cJzq9vGiw9JgSTZ5ffp/tueZ3TwyGgBqbplvR2O69QAffs+
4Dtz0Bp/8p9Xv7+QHxMzmItCpiCwPlf3e8DPlYOJszaiZ7XDDgajfaBfSKV0dalvhvYqO6ANl5Ta
kClBkNTsruz5zMLAuVKK+1N8lJ3I3WQvKNlLRC2faeM244krKY4+mit1ZR9mQlSmiFeQ87ipuZaD
Aez1xWMAwxDo8L96nxtZRlWzJLmHI0HAP/4nbaQiOV8sesAP/OLQTssBvemIQfslhkFNNO9StRVv
aVmYeqmVyIY1DJI58eSk/YNrLMYnu31T56Uxy6H+A7wXvfi3Y3aO3x8ptUcaW247JiLug45kLoB+
0JnIkPkLJ9MAo9puWM/Sw+ZEwvu3JQDzZvIuihRmCgL2I1cKa1Wmiu+yClSkLRPx13qK7y3pe1Cs
LIIb3C6NC/sgcVH/H6s+jTEmWcApbyLitePrlEsKXR1m/ve0GUMdkjTtKeuxDWaL3qJp00ERfzBG
ybzMelabQaMqpWUgh+VYsYJJG6dLD+WiqcUto0obHDpHa43EcKPhnIvG6VKTb1c/BYammhUn5/yi
L8JZG5A8ZcxZrn7migkwSwp/wEXp66scFk+Bqad0cya737kZwit4AXPR1DbTgRYkLXbtHNibX0tu
ZHlVPeh1ihLA9pdfFossFyBUlBjYZiOW+ZG7j83K0KozlJLmV+52A6/p22qgBpPeNOQsOGOgp82G
ZW4JjnUPtwkQ28pIg9WHWEwMrm6pLJHVG+wbsz8o9PLnfuZ/IUqQ5I4H8STo/ISHEB67hub41iIQ
HHMLf7qkm+ht8SB5MsvG08TUhr/xWkNXOBBDLA81R71vgo2Lg3nSlEA6fFM/+Tb9aNlFY1S/RfYx
fXYJ68uzjaFfuqwQn87O1cjKeHUXdTERsEiPSpd9ZzcA4xPjm5lzwgUyNz4II5ACgiCwwXI3Rp/G
GlNGpN+T1/p7j3gCjKi943ZbIuxTK8eA58kpyFItO+gIBnmYPFdiNnFNmyBZZKXAd1XfbBEyt1aT
6tXo8t6S3lUjPaJ4p3ApUl2T8hiE68DHDQ9DicVs47Hhu8E4p4543nDNMh6Y2rgF70eyXlmoIvRn
QRaGB9r1reb5mwTGmV7dRlmQQ7cUqu5I9DSm2legiu2fgHOazvDck2EPcyacwS1U9bMn5AFn5poj
HbXa7koJriiZGVtLtpLYstm/lOV7lrUVAZW9BLSC3VaidSDKYvAEJED0iCQrm9wWuf6v24AV+6/A
bcnJqGWYzRt+Xq7l5mD01YyxJUj33paHOX/qIJoDaOvhSTFZfTfgElzAuWVJsOLgIUCPjEl5pP67
/VmFcKGeYDgfuKcqBCO3klLGAIkPZtWBYbW9nZANWk+W3+Bx517v82I5KXI90PAckLwDaUlOSwKy
ZVBMoGAVIwlwTtonz/iHt79xsRQ3tfw8Sw/KfWsgS9OfJcsHQzvTdGaFhrIJVYlJ5yKA2QO/YGF4
tUVtbYc7CrquxGRKstzij16YevA/NHMv3O9zSoW8EIopWqPaR9l/K8N50Jil37BIDw0a1ikiRHKi
pexJ/Z7wO9cmgL2eTQXQBB9CqAwZRU5+pvfd/ajRNrTsFL9qUgHOqpcOYENtdGwJrOI/dJjfVZaF
PStZGlQZjUrIcXQW/7cOyIu0d8VyZfAnMevpJLqmfpW/ETSP5v1qO2TYCHFDYJITXx2nlD/+wJsR
kocgiW0e7tfIkbOPBGMujvyLuzHulW/KTMr6FfgpL/EvHG6pgBqZtMmYRgop6yY+6FFb6ryur8us
L8Vx8LH7oGG2PGPdSzKIznBBsD3XWn46CqrZSqgZPsvfkCTBA77WSRxcWZmkBRpXwnra2BXbspvX
kVLqf+aYpDlm07mxktQcR6z7Ceaovw003+DSFo7Ji6sxLMOX1QnwLf3FA2+ToS5htfE3lhsT14wd
XGKErCRoNEQzM8wX3fsRLQLlX5/0iA950wnvUDy58WTQKmSYQAwdAPB9kXbMYYUPEAbztsf6DgSI
kGUaD7qfd9Xh0xwqu+xCFERlcpgA5D2FD3fGdHOxe+0+PF0c2zDs/VjpGQvIooH3iLBx7FLO5Mfe
d+zdMifBulwa9lCiPU6xojmKT2w40i/RJTLcHZRxXh2XL9BkZPuCn7G4Bd1lyrEuqNDrOHyhcivn
kmXbvOzfMEYY22wsKulyuTi4fCPwDNeDiagQo7Zk6TPM03T5ET/gdpsitbcih08ReTm02bCJbVNS
kHRa+xgoe5njnbV6hu6nESvr9m1568N4ZBCAATqy+slhMjNxTE/o4355BYa5uAb/8r6mmH9Eoa0z
Fh5O3WqPLRwdgbRe66CFfoNUY8bKDU9/LWmZRRJ3/lK1iUbSIp7mt0SvY7amAZBjfoMQMhYdO0bM
9WnnAHuAZLZXsX+WMMJS9L3vIlqZS2XLMjazuMqctYhI5g5N4YP2XKBxskO0g8Z8vlpjavwJE69C
bZ3SNGQb58Wbw8TNZ7VAjA+2bnyjHnPHRvy3QWwlQ5DKvqzNCmJMIaWxiZjK8HkKAlZrEIzs8CDX
pfCRsxHy3lylrwadQ5jbJB6GLyj3kqwrjMRFI92Lnau+I06SugObfR8MrcA/4EMFDHfpro8O3Oan
TJOd0Y6O4Cq4dw8RXEnBlL12NqQ5ehVeTlxlfdrq+OvgsaLpepWh3SlPqunxhilLaUQ08HQDec8r
4fnbDFt9W639yk+jyEeRxVhkVBB62TRDwXGLQvLdvG9rs4D4Mp8POZGyQVURL/VPrL3IY3a4J3VQ
1WW154RPDFGCSypDXJbHtPpMeUYrkn9NJAP/x2J92iBxBekbug+gYst6ESgcpluJLXYKH8pM8n5e
AnckLwUNcjbo2Tm/go/ZWHoXbh1XG+QvtyInNWTeHyWEP+YOPgk11vTUwkGJvQdr7WDpsYTiPWi4
vegd+t3hX2pkCzTwhM/rIYFLRJJnyAFTeWziOeTIhfHaziAt9yr1SXNnoLHKxvoYCZe5q9+CDfMR
dLwQ+Vxl725QHW2ZX1orbNZ/6sBG1DlxFY+ehsMhZm9fvVSQ4P9MdyUY/CfthQQKgslQcrg36qAv
oxlffbUwQNcqz2mgbGdFIwQFWxTJ94jJ0ui2+l+JAyIc4p9xD3N6aU2D6+UnN0JUVFbD7Ptp5idl
47maQRWAgLSiEfaEqjXTe5yyCRffYWRdzj1Q244wDSWL/vTim624nWeIxtPpWdvCAgP31fXv03l2
PI9j9e8iSpbJPGW/6beKtysGkzmp2JVCjEXkNRaWz6R7rNfMBdO0tToCH81SIaRuRt+FYvrHpHHF
j66Qje7KROrVHC8kIecwY6jn8j5B6VkV0JSShbXDoD8wO0dao4un2drkxAYKjPprlJJGZ4GOdDmp
aYt9vZUkQH3ZTo+yRtIcjgZlGpklMVYQwoKZvh2G1j2Azrtprsp6B6M2EOl7yrdejIgub+Kh018I
YMcoxU91LvjVOQHUXpXWJlf6T1cvbW81RG+XS+z5BXmiRt/p0tIPV+iEL803xeQIkZGqIj/NJaTc
EQKtKmKBbGmigcAwXTGdF/2cyX+HcoJS7yVRF5uLwuGf9/pO3ek3D+wn4G5/hiwqpcZwPppZFNN3
RkJNpMTYftFpRMU2r8LYmhjeFtCNsE/C2yqAVBB4z2NCjQi/hbAUYeo7udWZCp4xDDRGEKvGwPL+
yTjzOSTsMEcfISLLySLzvYgTLPmkXiEDJdVmNBgPBJCvd6Ef6cZ5X45640nQE7QiTlvV/BRx55fq
Z/1D9Px+mO2RAHHgVVD9XjzlfQoAwq/fxCs362IsF7TdxPh4/S7Z2u7YTUaj9RFbej2smDEv8kWD
3vg4dLoJn1YaP4UM0PAob35Xs2R8NUQ5h1zPjcgCWO7+pg2JujpM9+he6/0WohO1JsSDJJr0r34x
s/7oRkTcaTrjYFebkbe8LJr1jXZgHFIOEYddVVl5lMiEiLyS0i7znDrsXfgwP3LmOBR9LoqEkJfG
+OcaoDHhkje5rRlmPU7WiSQ0CS8UtrImdUwVDheAn9dBIkN/k25hDb9N+kMc4fZWxezMUoI4S9YZ
D296eBtSmYvEJHhJJgawzmQoFQRvNQiVjTRAZgWOUYdQX1qaBdTlGig/h2DZITKpbDDIbnnOIMgT
8crmGnWZREM3FmBbZKWU70JkO3lZUnnM66kObHx63plU/tsAnjiVZuaO1oXrNLk9K/2o9IcLFpGe
W5Nrw6fx+sUKO4vr7Jab57NGNzbSzCScAINyQrVGa+l/Cn1AeZ2majuyOJ4gqLg8LN8Gv7WC2Mib
GWamBnxIm5ywSaqC8s6KS2HDvvEvnZOySs/7J9owWZ6PAkkn5Azl0Vzz+D3z4qNbrF///lBX2rNp
ZL8eFxDYE0Dc7mNP7Wd8eNKso5sDPMfZAvyxrx2SvrY+VaXB+Iwh5HdF1aWYxMWeqMoYMyC5tM0C
Z+bQNgkylaEya6ZrRLmYpF6kd8DHRbyN8A6L2OyNJe/PIjUnEd7PCK/Tl6+8twJoG95UKuYv2sP3
QHfgyhuTiYu2LcTwSxW18lM6MM+1ZJHr+VH5LLhJIvVBZ9d+UuwED/h5UAkW/UmVe8lLwUYF3nmr
nffSAdg5aBle4c81zHE36Gq8WlSRx9TPfAJrFL7fspFgEMlwsIwVCatfGx0MXW5BDeAwb+ud3Qbm
WORXOiT13WevFHLcha0tg5f6n0M/AcO1j7wq/eeIlroF4xGojDD0RagepdH+tzyikaK2xbDoOO4r
s4AD0ZHK5Keyo7eM76Ru2Dj8Z54jYixe9LVqosxlw1opAAgsarHg02MW3T8mYvmwhY5RzWV9rBO2
pc1S1KAtP9Z7bkxTOTKVQ2BYbK8mMbeB8MAbL15ExM54q2QAl25IUaBbuBrkqGfs31iYvHyDT/vz
6bhfI82LMkjWWNCOJexVofPyHYjIahfEWbMPPRKURmNMqVZeRLYjsM4Ix5yUukbVINIzFQBE6ocG
yaSZ58F2KF1Jg4UVpWkJMwNXQzGnPxyZcnpGUGQ3Zj844/5xzcjlKbKrnQp1gjNd8taeK1gOxjGV
fVpS1D93PUA/5jQL8ro8pI4SpasmILVzBSnYuLWgzN5otOlT/1SPkjP4JPvSaDVoFhPV1qi9qg7s
Kgle8swmhA23MAV36y17rsBIbK/L/f6nffnIA9z9fKAZDnfOZNEotqt0rtNd29b4huGpTtZVvOFJ
RVNB7JM2o9IA1Bt5hTKq0SZ9ywmmAuwDX8tc8KZvLvf79BbHGv/5lwifK7GS/t9sb9+lj+scZtR5
QIqXLrvWLo5N04Xi5ownbqwT5NnQ/wMJOUSZ7bZLN+l4Vygd42Wn4niJBpPjhlPwqO2vrnkZ+VSI
8VLORzCh104j/W3CbtBNOoAFeYv5zOx54Xm/gaWDIh2ThgSZYsDO0mZnPMK9SgzDADMDBgVcV4g9
zimTb1XS3wjTEOxCDn9YG+LpKAkemdAiuASbwbH6HtvDVCHtjo1qom7r/L1Ca8IeSryPMKg16Axa
eD7MPAE0Ij9MtVvXdL27WNoX2UMRfKniIoR/v6433+kWKD2lVuEfmqi8TQgI2KIYFJLaQA2NI6uC
Ktjlxxn1O1Rxl9ZcXh1UjF3jBkVX/o4Xlcfs9AuWSbeBT7SbH4Q2+CLgnurcia8R8su2h4Sp9JDT
iyULjubrbPUSfQlDLgLQFBiy23jMPk7F8ZeKwlQMIKp3FZMdD/Z6ZIif04Ybtu4E9BKW0Rs3g8DT
Memmt9ubUzhXpPJfdPjHgScOU5uBBvkzOeV19MpVP89YMQQWHI1EMWTRKceL4mLYZPvKyMntrzdk
t4KDtezZfOPIBpNnU4JyUAoxgRuk1UOHsW6moe3P7ZuvFWLIXBAe78mshLcT/zUIIuPZpG9jTe5C
eqI3GUyr/lC9wyCISt0DVK6inAFBVCMwbNfbj59Qj+26kKC1BdYzIuuZhqKwI2gKadFZc1HiOJww
Gr0e7T9VovVAYPFSQhfKt5WyoN1x+YhFVqYZB0lYrysUxk1sMuzlPCPx+hbitvw/IcR8YDvJu3aA
NCgVXB7EWBOm2W9osEdQRYSHzIErizghkObTn476ngiaOVi8ratFcIqBFXsK6Q7YSHWZNuUVpN94
wvxCh2a/VqPFgIAdpeISpWDkaOjja0tpNUwELVW/kVC5wnYwdElQNkOgJEDZuknV7XN/fwxlIh9o
PGzktYLVMh4LNYSNM5tNkBK0xlTBNx60c+rVgOcHb9/Opjv/bQaTgVARmZcdwvuMkxZ5IsSS57Uj
7RtNpC5RdSuFxH6Rlwc8cqb+JdK61kK5vCNvT8MUT9EgdM4Sp+ZZDBUs1/5UZ1/I0Ii4wOljfZC7
9M9JZbeerpgD4NLQ1o4MLhLqLhYRP46xvtKQ8qlBFA2/D3orrL8tZolBigQywk3szcMXkDZiUcaE
6+XR3Y3JjuaDFSxZvYcqCZkdl8X8djWY6RQf9dM+Jo5zpnGHjJgSZI3y2K2sgY4hXW8PEzW+1EPV
PEEiGbGJIl0rxYRdyuKDs1ASzaGbkXw7rIc39JzrbzPLHhS57II4hiWqlQCQKpWj8+XBNRni9x1y
WFKGju6XFOQIu+HdLyVFuPyrmC3VEQZvqPI7Zfn3qjo0P4OpcXVRPafO3R15NMLs+tpm4Cf16r6+
nkyPKuPIFwVJODtgZrLG/jgEosFR6F4m0lulDkvpC2EVCkvTFs4ofNJMDOMuAMsbek5mouzZVQid
Tsbau/IEatHx7ZHoCEYF8iJwP3pWNcz3BeZv95eJT7pa13KR6wsrbk6H5ypCFo+jtBKVPMF3dFOA
Oa/cNo+X+JcpuUh9dGWKSFv8vVmznaglOlFy6p3l9xzP7sfVYHZEC8MvP4+9cfFBU8utjrtX21WL
ejPiA0/Ia+MzHfEjFE4ovOw1xzCcO77kPfLL/Hq80k5E2vLJfdg5Z10AAGWZnYSDeT2TnOT39R0q
zorMhnBPsuCh6DV90o+IyoZ3jWSb0UTDnwqnLVZibLnRy4hkaHwy7iAK5B1hzxNbV4GZYyiSErZf
9fA5iW0GEsFXqBT6KlwuZYLgG+F2YFX7IBw5dT2VTDafECoZcwJFXKum/qjPg5slavHknp5VvDct
wBkDnnre5QPfiEJpEreOqlUS443VNcnKmlajylvliG2pKc3mCzezll2qiZOdTHNsTlW7WikbcvEt
f1kcXYMEj3JZeCM2f0XZww0aHQ69D4vI+NuQWqGpVTmbHCbZjHrjlszhdfGTmmrBeUuF3oxBWuMk
8M36udNEtNk3RzR/bho+G+FCryp27m3/rDKVps4tafQ/KnGcz7Amp5zyeun6vAKgHCMmPMJaoQAe
cM8sdqGAa0WfKPYt2u3um0MH7KN97Al8YOEK9GjDzRIE+jIH7XajB3r8qKYTMIqfud06L0Mj6E7R
rPCs6uNg+gnpWGN+4anieQFmmvmhaPOykqeJ2+VLJxKEYhekR08eKLn7xNb4yPhfQX+MZvezc39g
MFwIKfCJDUMVxzU6eKy00AbNSf5ZKfMtMAxk2cIejtvvDO3h2EEgUCqqQlri0r3JB572yIy9CN2l
ltkRUwnT/9f3wcn38+OARkL4nSBniBqVlPkN9Hsl6pE2OgYhOgcwsuJiR3McTc/GQ9lpinAx+jfl
TGHGd20iq8nIogiSd1vQh35onHq1N71bR2prZbA35Doa1ZrfobC2cIbyGOvF6rSqjrHRUWMHGtuW
GgVxbAZNl20jh5wXJ2cT4dP5xx2BYROmxQ3KUykk8ma3O5MmL2OEc8izkso8S+Z1EKZPHRUbNkJV
AL589Ww95zUlu5rEkrAr18K9jeyhCg2TiC5CfHIPJsP4ZVCNYSmIfspSM5uNaQv0+gTr3T5gPB/Q
hGZv7hxaPOz7jVJxIt3Dti5hXupbW38WT3AJzX9eiex0YE/NTLp5dotNa0qs+eGnLMZoMEvHhD4F
5MgZiUkFhlb2RJI0XaJ5HImWHvuh6bDFjHlSnYlB/LfTuO4ynu+aQyriZDe9dmBmySJ8wE7m4p01
FQ7WRFsloI7twRgiudbjQcrFBjCrVquoJj3WmEQDSfpFR3mJwcJeeSYPkKUKTCOJayriXKbVruBU
j8sUGVogkLK3l1SAR77ZZ6pyaCRw2krMXhi495Mh1A0ITzDWDgAkO/A/jeUtEfnS7PY24l9q0kuo
oGQf/3yl3hOJIBL23FlUUJdRlZMVhobSVl8d0lGAqO1wARRhHinSSxwDG/fsyUZJvNuymYzwbuZs
EhPyfJc54oh85oUmk2cxdtd0ZRVqhI6bfrDi0KAQHfVzj1BYgoPGye87FtFHP7e3LKnWTxKTVB4D
eS120UkTAaeLry6sxOIgvy56jgjq+NbHFQTCtZDeyrtu5KTleDfJmiWvqUItZpI/PM3wd+7KTxx/
0I7jN1KdjzGIGLd4EDckGrNhxTIF4ELlNwhb8g6jnsRhjv+PKMCQAB3x63FhJuw6NZcP65T19LPn
QS6B6qhfvJ8BRece8UuCv6QYz/yMRQxc0uyni6S3yB9NkEa3f+NZgG7hQq5fJOt9ZJrT4JR10MBl
Ue9qbNqynkGh8SnzQodNC1Baj9QzMFyJqWpzagV/22wstKANrOkPzQhOyLEUljyU9RtwHdyYbNSG
hD2OonCqpRC+mJJYALKgCqeqF3P7gomDM47CJkJnAC43vaM7llWU3+wsWeju1jzi+r/HBtC4UAr8
S2hOgoS9Qhmbyh1ynLIeSCzYPS/iZ944ngiies8F+QZ4PFN16zfg9JZ/m36lV9VR9Zlg5ZnQwBsE
/wzBUJvTwsZrl1R5IkReCdeZZErqwgt60oJl5oTr5a4Bb/RFA0sCX1DVUXOkSsGLRoer+Vc4OKVT
Q0ShMPbH9NLfBEgqJlvrS1Nt5qqkIpIVf5fj9C7C8SCR/rravipDpffsBH+WXWCd387KjzZyYS77
AfpxtJyGDqD7PTilwlgdeeeHWwfB1tkOQurft0GrPXit9KqRpxMwIovcQtlsf1fIBhD63CH67bhw
Yfd133gPqsDedElAPv1C2CuNh7hVXq92a2TsIAsQSEsIfKbzDd1U+2QCEeU7VXcRDLYrSBE2OLT8
Lc6KUt2aCnFy7I3pRYQo6yUZx2QrSjFkwGjfggaTkKY85EUz/V1sMCDyosG1F0W7N7p5fB8Pxh9j
O+9aWkEtmLbWDLLEv1FG6mPZgeyZPclPa2Mo1LPn7flvwqUM1qqyXHstAOc8wxSo77OdQUo836m3
3gj/5aFsqSCxCbS1/eY7UIkPa7RrgiR3hTiUE86HyW+BlQusiHQyfHDLxQlAmCpMc6r+cJ7+gdU/
bMXRXHa9L2r55ADvJ2qcMWUE7P4dWThfEVdVrnis+KFyM+KydWKYtZO8gZi2xNGpomOTFjWDwaYs
qi8/dupuh/7Xsg/X+QIVSIFkBmWDpsEPsFLx7ZglN1fJ6Q77YY/jFe2AD0mDwxQxXF78xNsxcX2a
Cmk87XOJ1f4mAG3ZzbgJIJvnWOpXMVYvBXvPx5m6TME2cUrz9HQiL5OfuoXMz5D0gcq4gNxSNNVI
AfEcOurooLBPzXwYbZCsO0ZBVpPiyLkKec9hJ3fO/PcWjQjhWk9Ix6S22VtbJMPIAwqjV/qGfR8m
eW+i0VpNY9SxyYdX0Y+oETfa7LQ9ceKcLQsjvU6JFeYUbpwITKtfyS/jEj0DO1i/P2oj+iQ3SHsB
ByvE68iZ5rXrAC9QRkEp4m0E33+ekUlHNE0rfg96F/7XXXVQ7m61Av5nZBPj1RzUVUAZOBOgZp+W
TVRl+acobdLi8SeQyah4bE5D+rRR+tcB/gYmJxOKD50+YBKgbO6Vr5/nUYokeYzlCBnVc31yYG+u
3fz/60HwMmzSff6HitUgVRVAu0pG9eOtX7CWl/9iI/NKC6KidvnU1wzBMTyylnfPGGXBDnPoMnEv
zK/wxbqMMk7k/PNogTP7LegPF8jYoEzzYm05eL2nclrvFbWhnyFj+pM8LZa6kdDGvpK3vtREYAyl
fQOWRucTs+YLnBDk7tOnMU3Qq+z0VC6pnYb4+KI2m4lH0Z98/isZE/aoM6zM4rheP15jukdvknjC
+uF9JT0qehpcwnBa4pxigkk1fDs54XypwSgQ41Y+pn8zHClp0rVu9PX0uZ/QWULGvgMrJ9JufM1N
4/S+v1xh5Dj+pvoTFq53tyzDsLzDGwf0zhdeqNctGl6r5VXkv7NrvCV0rzEZXkC+rGsI0sQd32ms
/CeUA/1TovxYpctmuXrGQSXzCQ5TinRFYr2pK+DWRdP/RHXpnAxC1PG4lWU+Xi6q5875CIWhfFI2
+FXxfgZao6IAKdZV4Yutfd2GmbTrl2YR9bqBBVQRY6CJFzNe1BjHUW3u/djkrwK8GO4eYL/1T4fb
b2iRB1+5arWpZ1NXg/fFpwstsc6uyU4zHR4cRd1Ev+Pz5aTljw8xxogyijyVKgRT6H2cDw6T86Jf
lsB3Wcjw1caEkGkZPW5ZP2kWQQalt9VtbfEUUKe8My33nwNRlYfiOzEgRq0RqptqioQJ+NCEGVW1
Nigkl/le94k7fAfXvASJhYwDLFUf+XfRBcoH5YplC0Lj18OyXnmEW+MJEpmgdxfoZTansNvqgQyp
8l4wEPgcS+hwVQTSNszdAu/Nr92lHl8vgtJNdKHH8WwnMaI1WvwOrFVqXpthNF1TOkNwAT4fkL7d
fG6bk1dvEDPTDfUH4mhddvcLFnWmy+EJQfaYeMqru+oa4V/Sr5UqER4NCSi23zocjUeI+G0JK12b
MwxYBsQEgonBuboe37UXkKlnFvr9ixZA0Q/I2ievtBCpz3TSI8PlGD/JuZJB7H4ShYu1t6MV6P0V
wgGl1vnd4dYu5ePvgMrdCrGP8f+QHPnFsU27OVzLClXFVWNeafDoBNwJuXLu3hW8Wd/vxXTeXftp
1LwcV3A/n6Y4tk5N8Hwvo3dMqCSpc/XsrhqxWC/nvTYvCQYpxMEJ7Qq16AJp6tjhU3ph0ItPpdDt
fIAzrLfK7GjKK1LmbvmabVQsp17VhlhgA7TIw5ELuLNHQ1UjfRkdl7/v+prFGxakTlD+Q/BY3RcX
dPJKgCZxmYlOyCGn+vbFNy6wSCQLnng2rNhkfyOGtzoejRHWqPeqntpWkaefbWfF+Dg+/xWf4sbL
fgBpkwGKG7M99O4j3kyEuLVqGEUlgW6xO+nAHe9UnOvPdXDpsLkS/x15GwEXVegN8D+pumw9EqK/
bQaGuU+xsBAZzxmsnRgyHVwyhgtApEhp841eZqJM6sIPlbzfvNU9RBaaLAxfnhBqANNDvV3ADXwd
rMrN9KKHXP9hPJa1jQ4jlIWLIR/2KW5APEtqsRzoPSNaEm2GMy1uW6rDQou92dwHhL7ewm9EwvK4
V5cLJvaTOb9Jr591SmU4UxqHfpwkQrlPbiP95KRn77kpwjERqAWhxe2OVs6NjTJLgguFm4Balc04
KwxJ3bwiEskl5gjSfwRtogGoD6w9xM0DINBrgjaslfUkwP3hRT7cNS5jKLknOVt4zSOFDprYK4DC
AXVrJCjMM4v2LD5VIHGlEe/NDajaYHpWTUG4zZ2Z8gu1hqqV3WCYhHS2zmLZ7eh+LAPeMhwKOKIb
URp8vKS0+V9HCmIqIuqd0eL1B1fpqQmsF3qtS+/Sh2R8zivbJahpyc26oMyqJOpQEVv12/XZ3sQ7
EOpNeCKF6jp+L2u3ShiBv9VqqckIPoYUJX1LuG9336XisZKAFdlVGQrb8AHfrazRqnediqnF/KDR
uV5tPyxyAEch1wK/J2+cManC1SIT4pJXXx0O20T5mAoxO1AaSmN1DEUvw6gS+TdLirRDKXk0TH8v
ynpvk3CoOdlMlsQDA7HslNJKkOFUYotuipzBnue9hMAcRI99p4CMIadDJ/CAtahdtItOZ/hDQV4x
ezY5yJ8s6lREESOlNBQmCHFkxzGhj0EikWCQq4YhcJUOv9z+8EeXVkCAzbzo/BKmGBT89pJnIBfl
AhJE2l+GN26JqEHD59xVjuIvTi4z14DydwhrqdvcNqDXxAQE99O2Mwji30arQUXxVuXxIUDnU0Tf
kKxxw3E0LUwYuocPDOBNTYgI1TEZvIDfMQ1UBw+2tZBRj0gZf4COn7rfZHvxkByVaUnx0rIWR5vN
hO+Ku48lnMd53whAMYnCYmVLWOb/8W/1XltLQjqoHgAkNwSjYfwLSgwxLqu6XfwnHc2uzGvXSA7Y
8FVzxBrlj72H1UUJX9qh4X5rfAISp4AtOEC6eos9Ue7LogkiCVX3aC8FLJ8WYv1dBrF7+asMG+sX
5iRQUoc6K8iOwLh3jTjCcC1sy/M+n5s90K75TupUvcKZPXZX/rGhtKPdstg6TpcuiaP0BqEFdcli
GiXquAlN0daepqJ0rkBwPBbEeQI0aHG2KPR2Hv+d217yzfBrAYXLhGFGv5SfnrbrSndH8vovRFkY
u1ePL4JjvRSeSz9Byqc4ZF9drXkX3qGEjKlsXaurRKQ01UtjwLEDXkw2FzfUev0RMPj0wjUjADY+
SD/PdcktwhwutMHvwxvtANNgLFOWh6P2q9UPbvsI2lPWxO1COPHbRhsCgjKZe29PNkLahv539Y9S
MDNDKho+rQuVzjbW38xckgoAnMg9X6HePtTs79C9zoe2+vsY+JeNEjns/wZbQ4At6be6XSPW0mYr
x4hgzf9ugkvssbR4FCw8vhel2Dlk6ZUDG90kSdfVka+t8UMqLJJv6TivpEuzBXGdxrT6TvGK6Tpw
0Fja1xSpITNiJVl4haeR5kFL9qzsRn0e0ngr9FI5vIHndy3sRIw8NdJqhlyeRVV+UaJMGjh35QuI
n1E1i6RFXHzebwzH8jLt3N04WrIX2u9jzFbKExdm+04+E3lrRb1s8Ru8Ra+36vf4rrooltN4mjWx
ZK+OQXgg9nxPhd4+Vdkl+pkA9MycGf1WbnVcSYf2yHps/KNZypEc62I24ZP/dA013k+JpK5T9XP6
pM6Whm49TvZYn9IucD+3ueSqI5F3Mlh+0S3SowsDrVBXSqUlaquYi0rCEd7E+q3/cTNO4a0/5PRm
SzoQvI8rLFhA4n4zQOZjewibHStWRN+XWNwouiePDynXREfH9r05QisyuQi+fEknnioLvLTWPQZA
VXd7zRbYxjY9tzxWEC5OTqLleiqxF0/NiJvlhB+Q5zjQBTbq4CLAvpR6IZBKX7fZkd2yM+QBHovY
wIulK5XVBn0+bChJdMkZW28Q2V6Zu2v6qlMCW6DnQoIU3al3di/3umFVepJzX4tgv3CGMR2QG8Xy
95YrAg3EVRZT/bt3+2OkLMEWjnZ9yuJ0S0vL66OX5ccP9gtpoKdlTO5nPxnDOijGJNemBTAzcp+J
hs2e64DJjW0O9qAZQFAj+U4zZZl388WBIrCGJZBipzSsQ8pjoS4uQs0J2xyrPFxQJj3WLyY0DIXJ
m7DZwPyJI1XAfe18T76CeNYxAGbnqpK9kUfW6Vw/PuJNPSsHQDrsne1GLIwOpRZiVv6m8Gthjcox
Sw9XJA2svOdjf0401NF3upAyME2ksmlPBA3Q4+90j6VZSTztC8lIaVwi6G/UBXUmGumU/o4eROY4
dP6UqjQRks20COWrm+G58NWe3wJ+0lROxN0EEzx5wiBmXaqY/BL3xqsKEYgWkxS0uXq4flbFDRAo
TPk+NgPLfBk1IOPiUBZjn6O9/sGd8ZrTI8REiQ69YUHCKx0gOI9FXvAeZCqawMBT0t7zYkmGQh4m
GSX58Be6odLqBtRZf6ZdXayov/V0XRcqjPmDEL2g6EW2BuyJ4wphNw9obZ76aO4NOx8IwR8GU+eQ
uEu7tnVI4GiW8PrV3EYsxZpaOKkN8INTTynQN2ZOAdQN41Jc0cL9jb3JhrT3+bi0yJ6wELVYDwgI
+iCYe87QRyYPwmoNdNC18kOKmvjpRMYodJDSYRPSKCu5o9yundaqBgRze3dadmD90XePZrKLoYlk
2XuxLLEPP7Bx2SZ+BqQD/99ueLo2UaxWvFSBnxY7qv2bs45JvbiDTPmRY5i+otmvySViE/Dnk8Os
6+h/XMZWhEqRwHkXhJJduzoSfFOPfOqT63mAehgpkfX1X+Z5xGp93z0r6Rr3PYFmqAg9sGHa7vHr
REOd9tBsnGaK0+UVaRwmkbhxUoP3Q3yzKAPKleZAK62BVSq4+u5MuhX6mVD4ToJ6RPXAnCTve6e6
n5mhjkeiozmAeHN3pjjOqx983BRVpayFOXplxSE2P6ADRtHbE5rOMNvlXh7mCEWI+ZQ9MhWix2aQ
sv55XUVtzirz7aWw/UrIk/fqKqem03iXbwuDR0+kFfrTib/oDyEoEY+ozBC+URgQc+tCXvzbpyI8
s3b4n3feph5+KNnNoThuMISXWNgZR7Sx9W+CMd9TwHteau6yHZdOqGL9++coaZchMloiMcnRRgQv
yW//j9hMbqCbxFXfpaZDL8RvH9c1ZsbUCA5cg8PaA4pXfKat0WW+TAlNmaT+pi4wLwJC1JpZ5hx4
XhBB6sZFb383nfKSSi+7mUQgtpfCsvHWnnTJMIQkuE0YHHlobibFjhLT+HN07woLMdI+e8C4DBN8
aRwgU6n0O/i5V5RxfITggdwTTNGVR27o+8ucXS5LYAck7rAb61+yf6i06MI0v1lg3E7FhPt6cSoM
csb7WvIAjXUxhr3UCScDRoSkNlcD2l+oKm7fpVnrz4rI4HAgcefRnc5Ky/gzRvRcNF11ctP3MGuh
ylJOlxOYxzEoJFv9JPvr83d6V97ngZieXwnLxfug8DMC9tVeh0rpr3IiHfVPRZs2WT8Qwb1P1qkw
83iAAoYm05rJdW8d7avkjAoN+dqhffyEzpHuO3GvXuF/YLdrmhlucLsBBRw6MzONpRh67NsB+EI+
AxPpt28N+aI0UBIS8mCMVEDBizv/nrEd+ATvqAfqm694UBlPyoGY384Ove/VFj6GuQoWF5qeN132
iXsoiwoapluHJKcSVwcYBJ4hj2qNpiM+d0Aiu/IT9KBCVeubyKaWmY6fHenMRsnH7h1+mc70QQb1
qPJfJoc2GVYQtClOm1G5B8K02iZ+Ri6JM3Bh3nWqgocAWFskgnpzJHpfUKWPlx/7Un0pR3710dlI
zkYX3WsYdwXzDrbzayDXKSymqnq5JYV5TXa8eykIp/Ijn2tjQZ5tavWV9nG/l+O6mD3iugx87MmQ
bnO58HNRdgVScuFrqP+3WY4OWT7hSn6grF31vDyVGPNnIGp/b04+Rr23dhvkWr9QByEMsePmSH+/
pa/S3TisWluxeV8caqOyCt1Zx7cutuIQKkLYgFE6EX/vJYjVLLOnWJ8el1a6q3AQm64HVE5oQePh
rNCzC5mh0QD4QrPxnVpXSm+8HClVaiKcQErrxe25I895QRuPNrTLksG1eVxQ2cdsSBzlnrMqdcZR
Vu+JdlapuZDrRSdGUxGQki+6HwOcZ6pag+80pT8xQvzDzylbqwAZdjZ+cPODQ1DeIVJiaiRtSTTF
9nHMVN8v29/p9XcQ28ZsRJBGuKXz+GPoaA+WRDAZKrbTwsgR/qzNiHtn0qktabfPIiLWhLiQrLFm
FuaWDk3prkudA3UhttovBc9DJSFgWSP/FaukL+h8YLghiTjSX145maK+TieTgGFz8C3ga6yOu3+O
UIU4lUI5iJMB8PDEjPfyRvoS4oXD5cnb2SbJb9S5lkJZICFhRtGNaz4ZF5kx6sxKJZfq8bcIXsGx
vo6yEJJgJD/y0H9n6CpqZIpUYfZS/Fjwr2d48xx0FBkFEoSdCFF4wbXTiJp3T2EBIEXjql+L9GZz
8U26QWZWYiXzwkkITKm2MveU1JGiaXWdfsXpplJqi4oBa9BzFezEjEHx8Hf3aRYOQ2XcR/+O9+ak
3sdtX7JeRxTOskpH1+LQf43RlkKkK545i375H1bYDB4/Z9cGLg6e5WfehSnQaikUgaWjLu7Zvj8b
Ipj6X3J6JHjPspq8ErWLYmDUEC/m/mUCh6CIw2Y96LHbY3/AUA0NMGHuVnikdKG17zA+I/czc3Xi
V9ZJTWvNAs6OnSCo/wAlDilt3iUmmzQdydU/y2XtxW+KI+2t9blIRWC0u3wJ3+PNAb18qAQZF+sD
qZYLM3VCu0aH4rjEIv/oKqwgRsQ3GFgp7gwwy8GjUgx4ccrucYkJSHqyS6EcOqma+9HZTSnNwPcj
wtoCUmEye2yTnaPQTkoVY4JKeGGAdw5BtuqgMUreA11e84JyMOKoi6NYxDJs9dvj97mrKr1VYPKo
XbPmbu2GU2wOOrWFSyVoUIfJmAgnO8A2aFf/a5nkBI52xDwLz8LWX1xE9kzPsRUADfTpaeEKhgjL
cv9hy3MqR7AdT48Y0G4JeLdStD5/k34Hrl6FCCsRgYB2k5v6RunGXyavWvBaYqQH/CxkLXigivjs
8FUQIuishjw2PhY8wZZP+TGMLni60rS+xCjNt/frwOIX6qk4ZCgsYQ80DeCLmTrWwy5EwHSffdjU
hXG2q9KyXhZv0Lej2po2zA8sGfsB3JKdNB6Xo41XCWRC9s6MAUvMGCwJGf0M3+J97slhXKD7EJ+D
C3OOUJXTP9QIRfYkNn3pyx2c87AICw0QNKQiBmhU8W+nwUyY2AioK0gQQxhRzTUhsMONtZkP766Y
toMEe8dvl15ypnMikbfM4HGAlNzrDkksn2PVxpROuP86vYnTdQ3rGmwisYdw6dTfWNW+MwXc3aUo
BKpoV6KF8N74npyyTmGZL9CwZr7mImK1T1q8U1IYtG2+xZ9UhKv3gN7dVr6+PyRfycgAsaZ60yWZ
T2lWhLv3A+WBcCAkKkWeOhNqZeSIdEXMeR5luHbTNn95xUvo3fzSxkVyZjpXGliHsLvYHDEOWzT6
S6QGhFinrmILpLsA3p9w8lLGPBdS3v2vPVCUgK92LjujBwWyLu5UJ+W50W+/QZFt1iQJ42yxsbEf
z9CKv7cqmrlvjLwcw3n193+wWHjT2fDMjQoM2LUqepsO8QNJt2ekw9kmFed1QnH0cS1jmGltjQx1
rQVZgrZO3d5rU4wkzE008HSr/QT7wRn5Z5V90uCKZY783ddJd9yybeDHPu8Hx442/FP7GDpKXwpF
gHL1SUBnEOhTQh0nRBgRaUBw25/6oLYb9zZtwFF2shd3q6jlFCqvS3IExFX76t6AR8yumAffpgrc
FvLFoLoEMkPyu6F1sa8HK2a11n4VpDuXzd72FW/BHHWXiwHIdINOAYQAfmfehMAV24cG94W9O1Rk
nZDxFup4L+Bp/ZaANM91SRbxMF4ltEpHx3nWtAV5ZE1dSyR2/T/5iFdwiQhc+5neHRuw2rLNK9f8
n6pkQ/E6r28P3/RiVu3NmR2ZNFXfrtsTaKp1rXvaZh39EtvXeG9JRAtk38i7IHrHenqYBGP3Uk4L
5hDvw6IK/6kUCqI0EL2aVwaE3cJOB4GbV87E+B5a1nO9JZzz+RphzxLJT1LcttSPpXkGe60uwjN8
elG/jOXMWf3eC0AZdbzAhZz9/hWw4QI6Ap2ef91oeO4/2QLTs+0QM7OG3t+y+abO1aBfFPYDe+xD
Ia6c2DlhkOhlGG+mddDxz/Mb1f6NPb7UwTt4XfzAALbv17iPZCSnDxKBhRcWUcqbMDFtTj+p3haE
n8kXhsDyr9NEdLUKjCD5+O6jQu2yv4Ew/TyqRTnpDsyuGdjCdqT3jT3NEDt1pgcaylsChcAu3VSI
TA7U8c6HKI3vyiK/McWSuGAtzUeI6v+2orYKNto5Rz0a8bzLN5IxKPGFVvgB9yZP1hy4764z9mSi
+Min7ndGHS+JdRR9DUZ4bulQHBmnNjfB672LAggvalvXu88CMtYpfKDwYnD5MLVamSdvjMPzsgn+
lBTTEVWwpiSj6rKehvA9nhKTIhRV+RrsJJW0NgM4emhONk2w+9wq5lQRY3MAWDCXt2QNU2/twWZH
3D0TcJqHPi55nJYRN63FAHmkbRX1Fy3OkQRxvFRAH8Uqf1msfQ8dBlGheVpPPCvLNwnWCaJyL5LV
vf93OlRRBuzd1l64zzZCNBXcLk6IHLfThjvc0IApuwVU+2JoXCqPYMhWOzUxC+K9tnBGzdC5Kp9H
YRgbC4sJg9UElSRVRXGzCN3jsbwR9+rOWQL4PLeFYADatw3HI7zkB6ujU8t1XscfMJX0c66ejKcs
UjNfJZtSfmGa+sYDT92FnZG1ekQdke7GeEQubHE0MtkPc+QOnXJ9yGfred8eWmNX3kigmFnYruwP
9Km2LBeZekenTpJCO/Zz1dvWe/teGuHTySJwC6qMZql0aIGays6HtEyEojTsOIKUOg2/4daVSJvW
Q9IsKr04Kfok7McqZD4u44WUHwPzHmYGayTh9hvqR0isueMQJSuiFZal4qDa0ZwWfgEAYcy0548E
BinLu8VGBVKfgwsihsk1ytq4xUf4R3cjvAbxqiniumO9w24NdJOxuRlA2QXd36TMCIbeSfkUVCY9
dKUgaXqF11S+FYkNC6cVUj+5ZUpbLfAi42K6uRVY7LIfDTxf0gbF1FXnZshQ0RApIyvMJ4hHWUDh
ujsptCITn4w/sKPlpmD4EdQ4HXHZKPADn6scaQQDChqswuIVIxRPiWab/xuDD5KaYrkhkRF3AaOF
8sls3ADX6DTh5ang2CYsCiHwE+G0vR5DFUGoXYmQjRZcZ1UV3qNyXXz4Sbhc7RG12QC3BwaCw8En
YrMS1oPJ7cLLq7xPI6SkQBYwOlYTv6qVfsymnCKpcsAUXIn1e5QQ+kb85cRDaklGywklsNIcNDII
uAQ4IW90G+TcXBUyhe12BPjIP6un5/ojMFfhdhH1Yblpx0RRypASArGHaUqWIW61i9kDgHOWRIJw
6o7A7huzKdaX2F9L3ddpq233s94fp/Sq2QN2AWcTDk+qM6PY2BISTz8Zt69Vef+dpVhOkLiQzeNH
8hgk/8qn9rsU1/jwuJ69dCxLyViJR89H/z4A+pLQHGjOK/rl0GGFB+IYIT+eTw0kI6AXnu/rWUMr
PgkS6W9ppAfjWsmrMA5UFDmw4EWokzXrBd7B7gJdUq8xfQJEARBE7wJbZQs4xyiXabg6axUw10T2
gl9gSk4l5QGfEIGkr8k3aCTnSXqcyyfAbvA6k9VLiBse+9znpg9eRCouzOaXPyvWm0V+B4bnPIHp
UO178qG/oO3eCXp5390nT6ffiIOouyeg/FQkUQKrWIfZuep8u/RAHkCxWaC3YFBKvycRibi/KCZL
ajw3JlgYHcq0hnzOp/6OgG8Cn2SmK6LAWrjIH3Zib+mPHUuNhX03sdWQyl/2/EtKDyAXRShGcvyZ
a1oMJTybnoE2GyAcFRU6w8425pddHG8CLyiO6E+OAwZaX6uJRWaznEa+HcJVK4sA8EJuZi6pJVtZ
J4aTeVEzLMac75RMZZv5xIX+RByQP2LF4QTRIR/wcRxBIZv/46czqPwswFkF6l1yn96LrrCRhVmr
WcikvlWBUAqo8jH1v8gV5FZUbecNcNo30NCbfSIZ/f5y0pPjxe81N85v4BxJXsm/BIC9T5OjRRlQ
vcW9SFSCllywRpE2/mxFIgwZ9ASue6RkRbbphZfRjEdUApCGQEbsO2yVRsvjLCh8092ymnspXueB
WvjBzOZQdPxEThE0Jdkt78GRfjzlllFjR+9GtOe23dNgEFjtMNYPF4HG0pJUAtU+Xjo03VVZlT5e
nteKCmB9O98IpxoYX9a6RaP2xW9tukyutOsonBca988eX5LtVZePh2Hul9g0gTmAvr6CsZtSGRlS
lqEXK3Fk8ivIJHfMKlowf+lt1dXvGJnAOEDuJXqhxkCPxEbt8urlsEoe+39iJrEpzcewrJMtB5Td
uzXK6XfqId0W/gfWqOmLYjGrGv1AaT5l8LQlA0/X6gBy6AlTg6VqHEucgeK27BJQLumZ4jTorS2P
VYIWpDQNzjH6ZJD7cskDmaCnmVVOz1tfimSAV4KLZTonS+e3R57Z3Srcdi8F+mrf9PKpKexF/qiB
QiPFFVGYVnzrLfiRbyIYgk70UlkWihOKSv2Xm6s5AGXtidGmt1u1CJMa2xGqJme1asP8M+pRXy3+
m+9QVEsB/orYs2YnlSMgnN2xZd9CnbBdKvVyjDsNMSvX/Uv/CRrPoGJMuh/Wd0Wm6tnO6zz1LS82
RaI+2u5VPxk8ZdWwD6g5ZYqgbcrpfKyeBKl1tn4WYXSt7ffj5gcGj8ODT3JAMYy1Jrvz11Y4IerF
7ui1Tt1I72uuOGRuXJHSZFx6kdpCJAlQXvnx3CspocYdT+ZNY62a3lWysJ5UlPVybpba30C2qalr
Yta+bf+IQoAxyjrTZi6zI8rmhU5QNTqg4KWQUESvQThngonLUUca+7aYRVDnDCxATZ6e4Fd0jZzD
WYoAz/J/q7hz2FoTrDNC6jsRK7vnseiNjI+V1M0LG7fGf5aIDewCcVNcGhuKhqrZi1h1fucrxDjW
CT9oEp55RYHo0K3AX2TmGgRi/9bhCYuaD7/XcPv85xwzjkqFluoAjnijiLp7n5+tJtvaNAWrTTRD
0nQV4iniTbuFI4gQMac0J4BhFkltM2wBqktARRgMB7Do8m5ZbIxl6kf2bWXyyRvln6oj85A7Jp8r
K5+axlQBLVliT8TMjSGMQFcDvB0sOFMswLF3SG3keqK2c/KIZSbOf3oMOxqYF3SOhF7UuqVTgAJr
K3BwG4wqm95UJobnw21+EMim6WDWrgsIrU8iZV3QAcqLqPwuFCqob+P6JWrdLMmHrUh4YRKpNF7m
o86M3xJeaEgmNxGxLWz/rA8n8y2yln3/jGUxeZmMoPk0v3pjnZ8cTXjxcxRuD6WJsay9Nk8OM9hM
z9Q/AmMlC5ZT6YwDuGkf8q87ksltRMWLecWHFGY9axJYJnHJdwcPZvshGVAfRLOUNYAypoXOy+54
we4owb9UHqSl2lACGPBGnxYffTfrOyCQ4OT9HEqjNXzUpiKbomdYDzszz7e2M6jouXF28u5QQBgo
dxiVJAXtD8pF4NvaVUYHeORwYQ1xh3fdLcn6DXFL/fcjH0LdfIrQdGYNBFDGb0HIuATuDBZARH2a
MFwL9P111csh2eDeWDYC6EGoKlbxoTUeE/bIIrQnhY7opNeBXASa6e84b1FSr6ibP+0wVY7lbUNm
nk7V3N9OZ3pa65etyd6CtfOtQrDXaokEi7GNzf2vWjBGmQbeyjkOQf4+X3l+UahDHeQiLPPkqwAm
vghKGKu+Is4fgCWCVTHo+tD6Rm0/ZA8SXtQh7qHCZmKFT6osEnWr21RkhTQ7JWBeYUVHNu0/KF/0
2MNUuVQuvuD3pegRy1dYkMzbKddRQr6j6+X7hb+mGl72hYMDez2HPh76nguZLbczrdwY9Aa/Z/x5
VrEVdki6DM4ie6iKjEeRtuHsu/q/9u2FPtavFD2u8EwjC215lPiFXkLlQfmwhrSMDo4ZqfIyb93p
zP2HE5YRMBRe4dHx3roCuqnw1kHFypOTUUJSSiLe95SSzAuV+L4QYkqA5vSuT/WVuOpVQG61NyW/
mCwbczxplLNofUifIOPaTJSgKw00YE/jsnEbqjACxYi9Xhwxhr6TzqY2hSDDmgpEyHFGAzIK0RDU
G2EF41aRXe2BvlOj87he0U248lV3ldOcErsybD+dohsShfH0mwHQBDsT+Fn7F/WOWCFTM0X4xaPk
J7SyPoRxm56g1Jb5n5EN0CDCMBlBCoL8hPepHUyALvrvHm95a9E4CvfybD0S0karJXtozbPGfdWA
C4J3dClhhF1DwMm9t+flz1L44DoJu5e/AqTQ95ZMUjYLYCQCwYeRww86p74BMId0r2TpsRt5h0CA
YVpV0wUyiY8ZVXJdQ594Lflde6EpXUd7UxnwggNeGXPwWbeQI0YHm/AhqgX1afNeUxRlOcZI+qF6
E/sRe1lB0V9qQbcRszU62z/oDIgfjniNuJBfhSS/h1AlZdqEhF/2ZsVEAxCTsrC4enMaXUy0sM1x
M9Vqky030NGu1MFfgXoJJPLvfrOUTOac22dpJ/zLUY8r2hK2jgGcrrHKps9oX/1jyE7gsIO+raTx
mg/fW0rFzdAXtnxglbAK4r0coKjoddNZyds220SssnknN7PVgb+vY65Z/ToFYpMIr3WkLDD4BLds
0Cy5jdH8kLnihiMvlzyKqtan7ZWNk7KxlRtdxU7WUcpSsarAjVKxGXUYhHTsfuRup2L3ZuKXHWAJ
5/T5BDh8yVMBeCzssC/COqDtmjr6PYDMeCj+cgWrws5LXKQi2UozYkc9glJWBewO0jgduwhr5Qeq
bewTA4UGaUPvrL/jOfWp49ihhCBq65gQOsD1+k1GsP2rn/ZPO5emhtGfUW3j3daAGyiVzEcqQRT3
NecSPBgP/sG1eQSwzZGfAXIKwUHJ/4PVv9Z5OT+L2lUkZgviFPcYQq5nPSFs21TS9AyE8xSGs/r4
yKmT1m165DSDDOGWXfSN5cQJuk/clKdTkFfeHAA5BB9tX2WXKXrHCyrsCe0+BlPVbrv+F9TjLGZu
dNFO0BLyNOlJrdJo9sQtrxGbC+NtSIU8fjtHkhnlCgRxpwJCgwQ1BcYh2hhpyT3zRcjnE4o9iaBZ
87gRaMhZBETebABXXgQXBgI/Sg9PA2ezxH+0ClZByHz/aKuaIRKVI4SFqDo9J74haJUpeOmozgfR
Yt+jo87kLlse09/PDxBOpu/LJCKluTIwET9jzavhC7H1o+jzL4zCjQ7UbLoEPd2OEdqEV/4goGiC
nOVdB61ChxjvuW/6Ht3+NBD8nqFtwAmb+Bxowr0AWoyFOVxxQBoI2+jSQYlxqptjNFOo2J6cdVU5
MQRwIe9GYStHJ8/7U+qtw+S+xsDZiP6vmw3ddYWi/yE8Q0f4DZhjEdtCZ972lsEFMk7zBxTBvJZf
UXTUPj5W8VQcBz6mEBjXnaMhz98V3RxZlXMeuf8VO3fv+Hkt/PhUtXTts/JjB/W1LWgqF8swv6Ei
FiyOr/y4ZKwWMwSvlcEXAp2T5/WM36Uj4SYiqgdi7uvBT50Z2x/7K78OHFm3Ptcl1GzZFj6E4xag
rqtDJxEjeYe+fFyyTx5EyezqJnirIKNPXycTJAXypWyjnmIznfDS9DQNtsegpyqVCEsjs99OdPBA
vTiR50rYxakLsKF5YmxKAd4m7AgfbL2CtS37Gg2eKRh5dH/SXQMaUnaXMapJvfXDlr6bI4rgxyzt
+NKxIALq4E9ESQTjZ2AaArDfS3EDYly5FNTussrwJnLy9c5mjwPfVuNsOg/IfsfNpeiMf8EXGcMA
2IGb0hsZJiFiEp1M2tByybH8ZBNlUxCpbyKez5aHFRjgmGLGqdvGVH0HQCzcxLMjZMB+I75esXVI
43TmAaW+6fm7ogLwZCfc8d6RgevttzHtPb6YWw5fNCrjWp2zWnd6Ozbk+AK/vdKyNNi5B9e/Z2fR
2VBAF74TLADQLzEBKSCCm0HXZO62Ml852AcMb73fE22NqCsflL+Tw3QNch7JEw/oVb0y3yca6ETH
pUKHrnO+KBC0hnzmkMEPo+HRQISpVjTZ9UpgEZGQ6IIt1lrtfz4b60FOIld0tFDATuctOTsJQRoW
xSAIm0/jV+XioWzN8awU2uGg8fio8hvv4FRk0hLJHjeGOpm5ZxV1pbGY7FTOXCL378sFtLxawanm
yUBcHbr2GqIvhp8mxqbXPTuX3FwS19atNAcFJRy8o1dKjj9hx7Ly+04NjyXN/LPYK0CFFCHJLuDZ
kEJQh3pc8wI767B4cPtazJ41IFqdy7S1qYyW8lf1fOH+/zs/KB4X1StodrKqdHL5lQO2pbfa6SXk
PcXtm6gAHJFsqg5Yz34OjTBbuuk0d8aNbmXFpjuEiRj/xM34yac7CI8DSG3EHFkxnt9W492ZJ7OW
rCubo2j1nFn4vwZmRu03ActKYzgVAIoQJaZgpV1X/Vft2dJWhZ7W1SQAV1SUckj36YGjeEJjhptj
H/WLT/XLvERA8iwKh+rA+V/KHqZ8W5YuqFsSPyyQv+IE0H6SBW7rc3XvILf2OfC/uBSobOTg0j5D
62r9Jvd8OsvGFN+4HKzwR9qptCYlp2wzYRQBa1xD8RH5+GviMOdE9HOZ7go82pYrrsa8TT63bxiY
A96qKJ1i6scfwkG3Jkv3wgd8hqXQzA/JNSEpQzFfdCUlukLrTfvDTcj4rVh+td3XWFDpN7omEzyR
3zcIy/DPBFdsahMPs+xXsRdXPELws3sXMlMDjY06tQScf//ka06vOutiuBZvchiGKtB6pYkXE1EU
qJcXwX3UMs0XZlcoef0YzcOenyOXaHYPYxwV3a/iHNv7MhpA34eKLrVy0XdmrK4ISMa8fOxyFqA4
GnVOsgn8RXAIHc1yFepAAh6rrtLHJrLmNmbjE3WinaE5ciBVOocEhUPxrPA17laR7i7wHylLMg44
46QzxxAMd/qvEOPZUli4CcdcBhLY8R4b29pJhKb/1vtSG1YWC+juQeKGUldt9omK6Erb+9zeQ7jU
Ts2vigesmNV+/RyoiPQPz/aSoDaTgWvPrQmM892wbxj2ZXn0y9dzwVn9LhpX/sneSx6xDi3UT/32
EPnuuFLC329dBmSv+tELKRwP6y7+Nojy9ERet1P6xOOEZLnxKhrcUi8WdSZ9eD+l01VGAL1hDH8x
5BGKzJaZxKPd9TZfONPf6gdq2vIO3R/evhT9sWXEtvRLHFdSMlkRoa5BTaXPBvokzCNaMUtT8J6u
wmCXXYGHil7coMDCVxVb5xSVjDbky5vf3dYEGM1S7n8JNImliyRxPFMDrXdKAPW40IKs0h/Y6+D+
BZjFlj1C1DlJ+gwzJS+lfu0E0O3y0LSNVVwKKofYgZsBo5GRu/6hIAX/cpMj0VFF/elmvN3zSFLb
CM/pf+bXLL5uaq5/Yr3V+bi9dWrYAdBHJmu8ewo9wsgMDgJeUzApZ38MbpTXoha93CV4z8k9XaHZ
JdSGknLenV1qnu4ZYkSfo+wYXe0ceOQVHLyiPP4mqraTHMUTPhnXPKkGRc4U1w1uwiWp02C4s2rA
h+Cxd+B0KC7mNw5TN5RIEN1reKvErgJKA3yR72fTrMlrN8KNW8nza3zC2Fio2FiPzIRns1b70tyy
T4vTG3nKM6R4CJR4Cpc7N7gaZ/9/+JGBSGJljrnTStN0B8BQa97CEMJZsrATe23gHSFgQzVjSoVZ
on5H17BpwWVKvAvnfauHsgVEw90HwhrRT4HW7zhiGGQccjTrFQEtlyFag8sxKQ8GpZe5u/CG95YZ
rWu5RYCW5jfAFDYtWPYsyx73gzXLWhRVTEfnKpt77VsUr5Hgli/5tvPaod3BVN0ucZrG8Mm4NVcD
Bq1ZjDjndzl37BeKQpbSsE48dYCG/QYX55AbRQHY/1oXkYyUxjKaU19Cy77jt+OeESIVv4owYdJk
kEus9wRU6UM2XhUeIw923ANKxsYEkNQL+tjvYFdJgNVvuPX0ZdP6VS24yXP2SDflvpFmHxBd2AkN
ao8HxQlhndrwGBwDFB7w37JAFPKqvUF1Owfj4jSwDDNGO0doSiSCmed0HPc6hgwg0CJfK1fIHPQz
V1dmVLAE2amacwWv8o7xa2KKpeSCHVtvC9fboMg26ZE8hq8LH8ZGsJbmbI+JCuNolax5zFNRaQdU
dXn/N8Baa546vhU3QWkzZQjObAtIEADBURp9vTJu5qIhZcqaunYbydMIqk/d03KCoUpYmD/q32cD
ZFW3ViP2L3zmIfaNpHhbrCYv51pwqf5WZuDhN0iT2WTYhN1gpXoGjAe5PdSEIzY7XS+byfTpCQGc
sqb3LI8a9tG4YbLV4ifb6M5wA8PRhi5JgS9DggpFJPeM1RQh9bYDWY6J82Zyd+wenagriaYguYsB
crct/9FOCL0tqJ6cvCsMEIN+9lF1XbBJFcWnXqnNi96m5omWKuVcgBl2j31X91uONyiG/25Begnf
wlvsLDYEZt1sd3peMMjYPAgoKhCLm9hFIQYA/y+I4h4Mae1+NBZqKv6PdqKcgYxcTXDdk1CdJSTK
jopcsgcsOxJQMbq9t6cwK98qXGrbPvuL4ozX098qlKikSOJC/fVTyjc+n/9U996xNvDI6xcM2xLq
0l90Yh2KsBIrZ6k3/vTMmL6SJE80lB6ihC4ZawzIHeucXi4LM7v3Wq1zPP4H7gq/JOYGoFFIs6cA
yxDiMNiLE5oZuhzpckM6agkN/uVq7CSf4jJ75vdRCprTwRSDBYxkUqus1wCFdVJpJCQ2x+Q9TyAW
9hITGS7aiG9gfxnCLQfJYylgirixmfS08vgoyzZHguGBttxC7vuEvjyXsFlj5W/ma1qluc8bpoca
mJdGkVQEhnB9dSc1U7qgFqBYpMX7ZpEKTIb8FX69Emd7JOsLdvZq6b7H0BsCcCy2DJoSUiD0Gj5I
lYp6MlDQDR+usu0JZ460ktWlOHyjr1gwXPyNSc87rZ2jhVsawPbaQ4q8YIfdXbaVg/Q70Wub3ibG
qJk5HkdBqrw0f/2R5j9MLNmnofmAVR/m+OjjqYKj/dyg/wk7UApF0s68pTL8w2D6JLtpAlpGDtjv
2RRcqc40nbR6rEwTiDlsO0FywCH3OoNiIikFyMeHSAOQG3xg8hW4AZkFvFYCWNW4umvLZtcFJDT0
dHsc0NFcV3SWH2xVaZuE+dbQBcnils9f3QwLvbu1IC0I0lnJzwhO+moCZ2JUJXxeoUX0eIPHfWIo
t7dMURtQzTduZkcATNsqAk4zILlPmzPvhOzutU7jXEKE9EWtZZQDVUJWAj2rTKzbcOTGcIpJO6xY
y2CnmQLYjJzlYOuzMmmlF2h5A0jdUh5R93rGpAfM/1o9Zd5qH26i0pETfa+zV401G0WLKaLseh1L
Ry53kscHU9w2Y+WuEi5eq47VeJWnXekusn/lWuSeHaKvWJIzlka17NAerS3eRwxcetdG7lVkNuy+
Hv7e4C4RIDU9efO3k1p3FTejqft4p4kQ5TqSbK9RV+yfyf8QkYyZP/8bmziy+Sj0Oeb2LbyOyKeE
KmpJ+aMvkbm7puXeVUvDPssvqNF/4/DrvIDfDK1opeNW3UaBmY9RxajiBFgthaR0g5PJo1HezHhC
Q6JawzgddAgnBwokYuJsV4gCVwgURNrgAO9iY8VwlRrrp6OJgEkr3Aik5GtGhbeqIL1jc02+O70N
N3oIZdM28c0pvahj2wMqUJakg+OMqGTSDbwlS5KWTwe5Tlh2B3BALsEr9zrq+CPbtWrJskcRhbdd
uYGIj8MhHlLRjg1JcqMhU1UKzNF80pxB+V6+TgtXZu0vMQYT1fXP7dfUI8VXr7ehZpzMuC/OeExi
xoJrvR51DDavfvJAwDwiKuBMcCqMVKOYv3d++o4gLtJNWNiwAEUrvAwivMypYA6cKADpBgKJXkyp
BV6rKs2HmfjhdKbK5yp1VfcPjgwfrqhaOJMTXtSN0iFE5Py3Z0OTLAheYbwWwDETHhNfepFEqJhf
WXELTHwlsTnlXqO/wtHvF1u/KMcV+gdWYJpeWswFFNM0hb037YNuAYVzdrmCAT79SGkoqIzalIi5
rd51gzKEVI1EUgrssQv24s1h3oEFhvBVQVd5uY3du0RjBC6gBxQTAxY6yMGl4THFgNZl50v5/Gxq
6XbO+EMvIny3/zPUMoxwRHeGihOzC+GrR3L0BjH9oWBG88rbphDNsxhd0dovPttEJfscn5DftjdA
ZU+DCETdD+dkbxczeNi20aqFWqj2CrWP0JDqBLgC+pMP936LNkBhEF+J3TLv4ShP+62+mFI42fcg
EvRa/b/JcLJ4QqWa+eIgqKNOEccERyJtGRZL3nly2t6B/AyTCEkgdCuq2dKzXBp5CQagGPZF/MSk
/VFuCHLE780yrAFInOJQlBEAPiMa9qPKPx2JSmRFADQSORo8v5bTXCfHCnOU5Z8WT79OKcF+O+GY
gLsQyvdBSzjn17QiOqPjnNp+Dd8DfxkBHLP18nwRrx+lc2P+puY1yAziHeOYxb0oWeIdj+Nsj6Ag
zVK02P5kHo53y3mOE+DEUDEgnN2CmjPDgei8CSTo3uW0iswyMWcNPiVG8+6txaAIoWREG3Zhtr7u
HUoD4z50zKD0/pvgtkobEmkM1lS5xRoqSBXtm0nnw3kvZBi2Cc1bGcmiWO4YKvxo9c8K9TEGKHzx
VGhn3qTG1YprNafyxJqon7mLeuwqluOyCohnMKlJE5VlDy6ok3jYj47cJqH+50GbVNzJqV8t+fbz
Dcs9WibN+ElXd601dbcPUSSPMzjByNUE+mF5VxTn3YRUAl1OOeO1RDbXQBk8CrhtXKJ2mH/UsSwQ
tMifMj+vQwUJ3RmzHjkprESegARUD9WiP7zcQWgRfa2o7eZGKNQNpr0v1287t2dfwt+Er+AYzmEg
9TgN9188dicMAXisU3EYt5EEhz+CKXR1vjQRcT+poxeV9ga8R6wGiUVoOKahL+GvG+vhsec4T6hm
3MIGUXSKqAca+tzoF1qr9QjpS4tVRPUzfl9KfOHQR+lFmAOzgsrtuN/rDTIf7jfPj2GWn1SuY0pJ
T28reNr0SUc8ln5xEbojdc98RlqMWT5ynSIAwdMBH2eaGn//O0nSb7tkBE6kNQj+2GuOvwyD/Um+
8T5Fe+mMHLJxy4Pl1PnxFnzyF70VmTWqni41CLy6MuKIGKELtEQPYPlqqoutNTX4AJC4ehcviOgV
9q1bRklcKpdtRtpGS33eeWMUOMLyYNTuT3FaGs3xQ9HUthFyUQd76RDsSTMUZFhSQak4LxoI+Odq
vs1HeCwH9ateLehMeWvTwCB/XybuHg1hrvfKTv395NDQBfOoqME864YQMZRHiKIvb81TfmFjY0cn
LC+QoYDUxW/6c3ONwi6tofVQFPxnE8ldPQT86Y8c8y0uh1L6XaC4BXJ9fVHZkWumO7CU8bUAJvxl
edTKSk+sj6WKPqk1v7vtSBRhch5H0HKmlVUt17fYO9ZP+qBozUQ3FO6GgQ8N7lB6ctFZy7CfzIUk
z1t6RsSv7w5+/9qbln7UCFV6wfs/zRrwTs6rw3PhmHilD9Q62FL8FrMMz/PhRSmtlTiOGyAuDLmJ
NTNTFP4n9jQB3iMl+pmvJddNdal4JCvIRITW8Dy7Glgwxur+8o/KJ4/O/A7sxRgGYNIQPQFTOSzX
GB2A8HN1Ef8AZERajJ6wQOX48r27+2QdZ5thMPF9lbfCU61EtJTXn3oIeMcktBv9WFsLDuNTQtko
KOo9fSOZpj/TbmvgVheub4rgL114q9X24AvI4h54XoiyxuaRwOdIEutNrlNj2Yy3qviAoiDhAYXX
d+opWn/ADbcv6jhRH2regJZG/M0gRW47wiRMana0u7CpOpduadOrXBf00Xkn8IWNtMCXDBKtLydJ
+eFPyjv9vVWn+4S+FmV5R9ZRiLRyZssgTxwujv0LkyEzR6le5XQaXQ+tRrBNTTw+Z3lVjt8XKs0T
K5Ykf34DkT4T4j5vjIEt1MsanaBB6vZElng/ZHud9B6kyFGuvgF6A2lWw52I1j/0iYRP5bnlXIxP
fx/ZyWJU8/RTsnqskUdfE9wSb3HsKlbrwLCEhwVWcZKCh+m8w0Hl9TCNHrAmRNlQhtwjVY9zmwU1
rjwyDMssmx5DRKxGt6QHDKoXiRvRxZmuYWN/XcnicDwBVTuwKZK3IFiN8suBimPCUsmi6F+YugUW
OYUPDq1JjhxOc1rvqohHot5ymZOZchWaCMb80qUfCPo+0gK//IxuRPAco/BnYMldbaEkf5rc3x0m
wuewQ5962FmB40Om4ibwBfOk/VNrXS7ncuwG79nGRDEleEuYB3tXYbPCY7wV6TnpaiA9lo212BmA
DvoSfalRcdpRHVHG7HqSeq+N8pyCK+ILIkQxmlQu/8S/5RaSN9mrT6QqliSgfzcfhwL1SB85E2ND
BExwzGL6F+0jww98C7UT0wKsbAtFiXv5IDUEh0TnqigJjMztheVIdihxNhCGoa5i+jMuzMTj4H0l
KdXrIXjPsn/mPAsyOrH5EM3RiUYdKXbhhXrkLzgT5YJG0uovayfAjEcFwhYYar8YFP1aRB8P6bM+
GVqOhvcyglxe6YDSBdi/iXA1Do/l4j5UF9hX/zEq3dLDbnwEapM0B9n4Eto9Sbw4eddvN4cYw+mW
bUoG1d86HDoI0H+xY87XX/wnE6QJwAGeQ8IN+BX2VFnHUWrodyx4ZbCvWTVCFSLsRc6TeJGbASxn
MCtSnRuezHqkdHB9AAWhwCiDS5K3lHhLhieEj3GljjkksKV6RpV2Gld6Ctl9VUoTxKkR04HQJl8y
Us1c+BRofWFj4ICvDuHRXsU8XjXfesI+CqM/UlcjhaDXmFH/76FP3WMH/49J8nFDfrPxiaU8HCWg
pYO27Yj2H6jdFGP4VMESE/9wssxRAzzRiWMC3piTnKI903Nq59bwOKQIhQbDBARC4wK+Oy2FZTbU
vFAWcQa9EhmD5Z/kFWY+SQQ8sBfOjAI1QAWN3ZYRaoLFiHBxlOmaalAUS3F3hlIpT16A237FOouC
JqIQ+4UNQK1vrqCVhCF8dykX0+ZuaH2VEOfafLssSVzkirmsCPZ6LIPLXaqm2dtWjEcM4Y6e3Ww6
+/DKNtLfQ+4j3fYNtB6VOvUytTt+ILXJ64+LsG7kKW+IymdoOZykCq59UltjrFLlVy248P/laEDX
s8c/VHGHYitd6tH5l25tL+4OsvgTKDuiUEJhlnoTxnoik0x+lkiwNE4sBWC+3NKGJZfgTc7jQHrV
fIiIJ+ALT8yt/lN9Ysm+h5lJu7A6GjNRDICA7qkFsehOcpCy7tlLv0TIjkC1BG3GpY+sZELYvoI/
WbjL/bgvc5tLo3aI7gJtqHGsPjpq8iBpfXRWVczXncNTfNOCRKJ5X2rJWGXKUeu7Qi0Lq/ugijCx
+QJECFms2ER6AchbgNpW3RMtMmVmFZK4lYl3uKHvJhrpPV1XL7i0q88jXSIq3TJf9tKp6dKTf/NK
dWKhYICZ2VNwhAxg5GHV66SQPNa1O5eyjvT9Q3j0Bq/yqhl4cpz9+Zo3AKmkO4cPEn4tQeokzBLn
0Q1l7S/wAib5sNSrVcLATKAW9JRxsHxZ7NNSjjeRX7HAZhCRhvUdiTURc1EllC7d+pSDmUHX2ZpB
/ZSBqJI3HnPpqyolqxx0CqwpJ8d0c3h6FkmPmj+i/Qu/EahtMovCRjPVmaK0Gj+38T57UM+ef5h4
L6rXysvwtVBP2HdXOQ/K1sZmfq1aYr3k+6hwyZPf0g1XV5m7UCZAIeglj0DDL9N3L2/XjUqA25x5
5Nwnvuv5kj6Jos5m53kpX9I4sxh/qwF6KCIPQRyWWEmirpZuMIc3I4DIfUnY69Lxv+3cMSiZQ4QE
H2+2QusuCxhsYXGcYJx9fn8KRmLPoy0GJ1Zk5R+fYw2iuJZ/cDWFRINwpG2YqVWUjUvmj4dBaN4k
AvuO0bkhF/l1Ebgho2Wv5Cm0Q7S7nasSyzHdFUkiNo8TdptnCSYpO+7LmI8618rL/suDucHhLBNc
TBfktSVAcnJhTWoLwFTx+jPgm3tN/ZAET8ku06HYzG3MYWfs8oKg5kfCw0655O+br3QSYnBjWYHE
cO2+fkR0mEpKnaYc/2wxP+n+RVmAjtp59EQiV04QWJpXe1pbXeSbo50uGvr/fei9qdl+MVpG3WVN
SWbtic/pcEXz4ZRjPyTdjWLAgWt0TZBavFFNN2WHUELSWSHh8nkkO/jY3HZiyKb9kyIjJZdVwRGh
PyqD5SFC7c19Ul+S1ZwJiRH1R35Pb9ZLVoCC9exxf80WKtt8GwJKZcpPamVFAW1aCnFLGlpzSsYu
Ly06rtA7Rr9Aorn+15pWESZ77ToMaxIhh/dzonmiEsy5Cz9RSSkCdAQKeNdByz8eza3Qw57yWu/0
5XrI2W4z8LqPR+nIe1ccMfxeCIP3UruxXfbo6fZHuS2iSlS4mIeDNo3qbzLnPUq6Bf/uGDAShdFG
7Oc1LhzgveHreQ6p0PB3AsffvdPxiiWSiWX1wrxsfptymGgVwUmcvoXfLDYWfEBoTTDENaK/FeAT
00gKv4BMMMU8gcJD5F8lBLSGDNikq1liH4o7aBD/IXaCwpWmmI2jswceUx00cSgBozXewg2ZjLem
K10aDrUzve5UpoaeThvf+4d3KYE6hQ+tHWlgMKj1lSvtYqMF+IU/MRRUNKuHJBlSY8lf9a7feyy8
KxSwBSjhidFHSdJkxpkHbSXSwK0rM7/kQgm7TlEyFGb0E2xlQffWcW3gJRdiYeFMO3h+9HK77dBW
9fKxnCuMzk0A0oqPxmkm+4ZuWnMIXgkAqnz5bnVvUBnowHmHJlSkSu7jg0a4Paf2YJIgkIkjxSHO
We/qJNM1DpsfsDhfEqUrQeyD0xN/M6+X0y5PEBnRzmKfqjCp9eN3mnvy//wzaLoq/7UPEba/Lnnr
rxopub10sb8jRy7YDlAIuMSlACzDKGpQfd7T8oLq6eGvOJZiKd9kZKojY7i+vZjkQaMQ1cbavqPz
wgpogC2lcwB4ygKT/pYOKD/i1eYJ+PSECbGL0cuqQL03/DN7x9vOk4793euP0jDVwx6IM7bp08ku
cFnHuEgzXFMG16hLxaNcMx2r6Nmh+ISlK5n0xa1zcVTLpMc9tNfViO/QLyKoTaRdDLUaWIlDHrAi
Gt2/VLsbK78taqWdPMvNZGdjLQ/Nvhs0I4T1me00+jLp0+qWLcTqrkfPpNrqiMmJREl7z/kfOa6M
eU/LiO50Dr/KdeT22bsT302wtzf4MHleejdhmki0+tDBOcLJVEWyWuU0wdoaT7JVa2v5pNtvkSho
2DxvTk5SHeVvFq6KlAceR4kMUsgvHc7pGBTtBHglo2uqgOgj0KTOpQZ3axElhEzVyEu3y8eJRAHi
HSjAAnqdBB323YSZasJ2OiLGciE9wrSTxbI4BuHFJXIT908zAba5pqhs6U95Bpl3tVgaE/pJVm4c
+v2gPg9Qj9qKaD+CzGRgxV2LbUZRzA30lAgD4o99Mp+cEL4287FR9fgsFil2aBmBMOeKTIDox6OS
NGup3druiUqRK4E8+kX8zXUf6+qnsL7lguuqCgc6+kAwgsd0uNgsHmiqgLPG/JgOeEIpI4AwryY4
t5Ox7SwHYJZ7l0Ga46aE6UyWaGgMpZx/RPA02fHKxx4BWwvOP+tTykmJveH2LXZsB/+5byU9E4je
18BrVJipQg21h6+7o5qK+j2NAYKks8tzxJ602TpRRnfoolZPbLXUCzdxW1k10PlR9PJxF50mN0dW
OxO0CtwKA9EeaYomOjHpB5rRoEVSFQSTTKlXR4iqA0KImZ7o0pBTNINU1lw/Lc4/QvhrCe/gLE0+
oCnp+7EPxHf1ICTyEBEHhtToWXvo/n0PdVv1vVx2At211MC1Me4ry01Mow3ZBeaZnVGD8X/CeSFq
VrJdl0oyqkvVYVoX5P/A7bNRgzBF30cRBJ8T8E9EesrY/HQvY1XRBIzw9dVPX4kDdYI5ZftTjVAq
fNgl/yETE09uK+xJQe9qCHnCt5YfnSoy5pDFglph9gyZDlLDIfyOmqOguS2dM3zkevZ9wHYtOy24
dbw38oAVvjGbHS6WsgHJQ4DGkSZGa/LwSEabNFsZ2sX4D3ZFzRL0kwL8Lox5lNhxMxRHEfua27L6
WmgKu3tzCU09jUKzs/M9OlTuEjwE+5iTVzc1anc7QQpkSLB3x9y5JKNTec1Ud8Vajp5uu0tM6jnA
GnUqQMIBEzNwuKOoLjYmDRDiLKvBdUtSISn/RT8JFpdJLd0rMn9WvRs8F0y8hPG87t+p2Sj8RM1l
xUaPOCnMOVBnXhP43BCNvAMvY7YgiGMaylSlAb9KWrQ3KOEueDIh8e1FPQl/5Vz7tj2l7DuyqZWS
DqF9tRdId04o2opwl33XU4vver3clEIgxee73j9encTpncZ4UbpyQcoQIN8txCebYdsxHmdnlxdR
HXI/bEDeOvD4tnVf46ndXRSTvgSdpDCOLZ/fcS8MXSlXZDAAKOwXH+6iFR7fgI62HcMEdoBwU1Do
Ab53IwWkvt2liIU35RsaFnZuIeU8dUMY6MMTeIiFyqHgT5OAJNo2w5csqxwvtJ7ZAKV/zPzwEjh3
3jU1YtppBdEKFSp0j6PhPuJiTkrTDLel+Go+VbXG24n10Z95/vWgvVOOb9URFsxcMYYZNzXifvza
puzkm2liEzsFCdnjzoHoEFcF5kgu6gZjrl86jdC8ETHT8phLY9HCPxVkMJ2v+p7L9QrCNZNnRRS4
Ncok5N/g3qhjRMLW7V4zZqP22LIi1eTm9PKXWWBTS4XMqoFOCYAYysZXBpSqHZ3bTz/8jZ69MyRc
lk5Mq5zs9qbclQDP2IpnG7QFu15qpoJmFTep8290uZ5q4g8Nfrb5a0VAri/6MTKRdZ9pHYOKeNcF
rvLbnUApm7082xsqKL+M/zklA3gGFYPH0xM36VfBULajJO8QZu6MtLiwVGHbww1AX+3KIjrq/DYJ
tAmMfbM1or2j+dkkZk5v0/zoDn9zCkc8wymJec97oXAS+xO4gk94NiuAnrZDWZQ11L/q0BhR3eUm
/Lth/l0oKYT3W/ZIBuFcYqEfWELAE5VmMWp/YdSgjTXN6bE37QWmU1M1oS4kfJ0+9x117ELoJaKK
CaKPxcSSluoLqdNs0htVZYXoY60TwhP98yfiO8TqiP9yFUebpRp0NUK9lFzinUudOdWagmQjtRFl
sdkMnOQOASrF/CNGeUwKgjuDm5BUFL7GnpI4W8xugpdMIfsbmlHrSJGh7x7JAhjwv6ntXQlVchZn
C4zmbx5fuBRggXxY3oVsm5eULnbo/cZyLYG3y+8Qv/9ANy+sTbz7re76r/x0qN8kKqvVRKTxaNaM
dqUZk5DxRytY2aFRhJLST6Td7Z/exayVpYjH4AP3ChagjED8y862yf931fqvfKlKYwu0lUQW9BUk
gO+/vtWVQcaGZ6U4ABGzAo1mxyeutQdjiNZkfO02MGKUMHQohhwsG5Yb1BA0Jn3DVjO9vfTOnEFK
pUuA+hu72/4hUF9kjZPPg639mGHyN1+PXbPLpxCs2PvmKdVNV1FQsxHBNIndzFvvEVyEkjfZBua5
DUJhdRGF6qjEaWzG8DTOeTULNnPebN08i4Bk7M/RUSYxeq07TIW80MgBww74ExY5L3ZAe5HxH+2O
SpHd6gFDRetrod20tFOW1dcUI4PGlsCQLEisPxFlfkMJ7byjReq2TLK9Wf7bvqtwig8odrp1hVWM
uZHxHfE6sZrMYkjuddKCYnVeGZR1dJmpuCbvGXHLN01KKHkJt2TXa6zCWRLpjgAYWasuCM3IHApv
UTXakMDUjjiPW09LJ1bG8e//SfvwDpuBuyali3DRJUlyM8N2E3L4RHd7nFnLkb2bW54YNi/yK9Ve
pMAXPs87uDSSaAPxc/gPhMAvQ6pk7fLCBIOTVAMXU2e6Hyl4ZFB5D2ZVzOmyd5vBx7HUJraNWNyO
Rgwq1G1oeF/cPmZtuyawItR58gVNVFajwEgcJEzuik/RT82ZBc2TBC3kclvaR85G3UXC2/efv/7P
uO+B2boq7XKk70BUc2+wmIz5A1YV8igOVrPrZQHRwL+CDBkvLEI0jvXoeM7qYobs5nif9t/UhkvL
Yl+Wq82bcPhu9b80Zgr9T04vASpMoAEK+Y5t6VWsiW5hbecOTw1mGpihKLSxmN+//mMYEPrfgiUQ
vTGqgitQfqoJ7uYLPPFEonjZ6efBIUQK7yTqOBfBXNkuXg+wSJ5njukuNa/xrv2IfOCN03ClmF2d
kGLzUKasB7FaS2gQwULUwTp24EXe7GqUSE8J9aocZCe0pPrfHjjZ4nUYO1d2TOJSZODn/J5NbR1y
UkzSTd+HYYszx6aPXq2Y2gOuOXQa6F+qM9ouVrzoZduHT4B4VvnNfQ/rF9w/Rtv6PZfVWj1lz4u0
ngkc6rrDhGXYncjPYUfBU6qFIvN3UM0BLtF1VCEBxIfNa+Y8X9bVRWULXmVfYldB71HWNmMCx84X
n6GsAyEl9Z9i9JZ+wCh0uYCKVeH56g0zqcsMt3QuU2GsmkpbML1Gbg17rT3fJf7/362Cua7zkELr
iZnRL3Ug6ElnpcYqp0yVVrHL48l14wEntwFrJGqxPcfcwQHNCmeQUzwtQGZ+1qFo4X36z8ZNbGMh
wQXlMzcMD912cxs7E2i0IQWxvD22SbOs1HE9wapSD80nFtKShNS5VyfVF/nA/kIudYbpM0/24Aig
EYx2U9BgYTMa+RekoByVmlAPWFliKx1FozQwkCs4pmlJskxtiRip089tak7enEUm3DZ5u1DTJf20
8ESTCli3tBO3qvNMAY2H/Bk3uA7hcDpuRjcWFO/pu6pDcriLDVaNAwdy0SL1ZVbeFOyFu6c+s1Tt
8MZ50bZINhb73qMdCfh6F1OO/GWqTZys0AsUY6dwkTyEMsw+bu0yeG0iFXvKnqDYBroqK/ZtJX70
PW8SD8fOFCbwMKgaMwDDrnJS4caeVpscP9HTBCTOn5T58IANIWNVa6joZEgZy7ddFUBywE1b2RQ8
VK/o43M1PZzyzw+Usak+PipuNX/N5MniBIp8nFdCXEgwVWD/5vhK2kQDGDbel532TiGr9V15i0Xd
1Ts9oOw79hDU2d48bKzIv/ua4SpFOpQzcOEukYJMUOGv+rsGOXE+n4IM4UDK+hOXaxXH5+mqqyWQ
y1yjfaab4yezbLL8TQ79xTKN0Ov0lMrOmkeW4xLw41eRvfWKFuAcF9zeGpjmd7N7FdIuRLyjUXSk
tf7+V+jOHvc+8z6oXF8nAEG5ko+cAsXvmCUxuoEU7uPMrZ5pjw1h7oEMHQW1NNpPXqE+QDeLc3oW
aIt9gfKwTM5EXaISRbKZuB+Uo3pQ4LXRPov625deeWdY8JrW0AuSeTNuWyn3ri0t5fGvpLCLjDdH
QVWPcsljNLWeP2vyp0lknZcmPKPn3iL5sjzqBXs4IB7lQ1S0zjs/URfXFhmn3qX0Xz3GaB+LgeTv
PRPw34uF32zi+aNnKiDnljFVdJKQ4rbA6Ux1vqTCCNmW2QqNelE19f9cKHggVW4ckjZpRPSkcbZq
qS2JYevt1O7hPOoL3NfX82i0iyxj9u6TrtveKaAbJ7pXn52FN6rqGuaY/OpBV/DhDf/ycvPHEjp4
OhG03UIPU9ptn4KfuIHl7023HWGxY4D8mlv4hCxj0Dd9rGC579uP3TzgDNJLaLVsaidPTk9t+h9H
jE3erLyscsuY5dSVXbxIXB62mLkqox6k7g4C16JwLbyIT6NwNmBEZRyQFANOBcV6/6NqY/ynNtYb
D5fIaGjv3h1oIBzvPImu4jKg8TSDXWe6NvNlY/QVNsU/gQPiKJwn6enGi05FqTkI1n31thjpqOKI
BoKBJ1bGqG0/lkYr8hgKDHmNRjHTjYwls3q4alzcuLb8X4bBzQjDa30vsJsB5ki9I5Nxopw342+J
rA0EW7w8gYV0xCLRHOJr2H52W4b1DD26Bb8hlw/KZrCf93WuToANoqkr5/owiaOQSvwL4kkbWiuj
wYuCZyAIZcCiyC1x+UlahRMdRb0oKEkKEzxGeafQrbj9SmshRU0ff5XqlQq1wiYD4R3K97qAvpm1
JBG7Tw==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw5a;
use gw5a.components.all;

entity fifo_16x8192_256x512 is
port(
  Data :  in std_logic_vector(15 downto 0);
  Reset :  in std_logic;
  WrClk :  in std_logic;
  RdClk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Rnum :  out std_logic_vector(9 downto 0);
  Almost_Empty :  out std_logic;
  Q :  out std_logic_vector(255 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end fifo_16x8192_256x512;
architecture beh of fifo_16x8192_256x512 is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo.fifo_16x8192_256x512\
port(
  GND_0: in std_logic;
  Reset: in std_logic;
  VCC_0: in std_logic;
  RdClk: in std_logic;
  WrClk: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(15 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Almost_Empty: out std_logic;
  Rnum : out std_logic_vector(9 downto 0);
  Q : out std_logic_vector(255 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_inst: \~fifo.fifo_16x8192_256x512\
port map(
  GND_0 => GND_0,
  Reset => Reset,
  VCC_0 => VCC_0,
  RdClk => RdClk,
  WrClk => WrClk,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(15 downto 0) => Data(15 downto 0),
  Empty => NN,
  Full => NN_0,
  Almost_Empty => Almost_Empty,
  Rnum(9 downto 0) => Rnum(9 downto 0),
  Q(255 downto 0) => Q(255 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
