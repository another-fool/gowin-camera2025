//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW5AST-LV138FPG676AES
//Device: GW5AST-138
//Device Version: B
//Created Time: Thu Oct 30 12:45:37 2025

module Gowin_SDPB (dout, clka, cea, clkb, ceb, oce, reset, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input clkb;
input ceb;
input oce;
input reset;
input [16:0] ada;
input [15:0] din;
input [16:0] adb;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire lut_f_64;
wire lut_f_65;
wire lut_f_66;
wire lut_f_67;
wire lut_f_68;
wire lut_f_69;
wire lut_f_70;
wire lut_f_71;
wire lut_f_72;
wire lut_f_73;
wire lut_f_74;
wire lut_f_75;
wire lut_f_76;
wire lut_f_77;
wire lut_f_78;
wire lut_f_79;
wire lut_f_80;
wire lut_f_81;
wire lut_f_82;
wire lut_f_83;
wire lut_f_84;
wire lut_f_85;
wire lut_f_86;
wire lut_f_87;
wire lut_f_88;
wire lut_f_89;
wire lut_f_90;
wire lut_f_91;
wire lut_f_92;
wire lut_f_93;
wire lut_f_94;
wire lut_f_95;
wire lut_f_96;
wire lut_f_97;
wire lut_f_98;
wire lut_f_99;
wire lut_f_100;
wire lut_f_101;
wire lut_f_102;
wire lut_f_103;
wire lut_f_104;
wire lut_f_105;
wire lut_f_106;
wire lut_f_107;
wire lut_f_108;
wire lut_f_109;
wire lut_f_110;
wire lut_f_111;
wire lut_f_112;
wire lut_f_113;
wire lut_f_114;
wire lut_f_115;
wire lut_f_116;
wire lut_f_117;
wire [26:0] sdpx9b_inst_0_dout_w;
wire [8:0] sdpx9b_inst_0_dout;
wire [26:0] sdpx9b_inst_1_dout_w;
wire [8:0] sdpx9b_inst_1_dout;
wire [26:0] sdpx9b_inst_2_dout_w;
wire [8:0] sdpx9b_inst_2_dout;
wire [26:0] sdpx9b_inst_3_dout_w;
wire [8:0] sdpx9b_inst_3_dout;
wire [26:0] sdpx9b_inst_4_dout_w;
wire [8:0] sdpx9b_inst_4_dout;
wire [26:0] sdpx9b_inst_5_dout_w;
wire [8:0] sdpx9b_inst_5_dout;
wire [26:0] sdpx9b_inst_6_dout_w;
wire [8:0] sdpx9b_inst_6_dout;
wire [26:0] sdpx9b_inst_7_dout_w;
wire [8:0] sdpx9b_inst_7_dout;
wire [26:0] sdpx9b_inst_8_dout_w;
wire [8:0] sdpx9b_inst_8_dout;
wire [26:0] sdpx9b_inst_9_dout_w;
wire [8:0] sdpx9b_inst_9_dout;
wire [26:0] sdpx9b_inst_10_dout_w;
wire [8:0] sdpx9b_inst_10_dout;
wire [26:0] sdpx9b_inst_11_dout_w;
wire [8:0] sdpx9b_inst_11_dout;
wire [26:0] sdpx9b_inst_12_dout_w;
wire [8:0] sdpx9b_inst_12_dout;
wire [26:0] sdpx9b_inst_13_dout_w;
wire [8:0] sdpx9b_inst_13_dout;
wire [26:0] sdpx9b_inst_14_dout_w;
wire [8:0] sdpx9b_inst_14_dout;
wire [26:0] sdpx9b_inst_15_dout_w;
wire [8:0] sdpx9b_inst_15_dout;
wire [26:0] sdpx9b_inst_16_dout_w;
wire [8:0] sdpx9b_inst_16_dout;
wire [26:0] sdpx9b_inst_17_dout_w;
wire [8:0] sdpx9b_inst_17_dout;
wire [26:0] sdpx9b_inst_18_dout_w;
wire [8:0] sdpx9b_inst_18_dout;
wire [26:0] sdpx9b_inst_19_dout_w;
wire [8:0] sdpx9b_inst_19_dout;
wire [26:0] sdpx9b_inst_20_dout_w;
wire [8:0] sdpx9b_inst_20_dout;
wire [26:0] sdpx9b_inst_21_dout_w;
wire [8:0] sdpx9b_inst_21_dout;
wire [26:0] sdpx9b_inst_22_dout_w;
wire [8:0] sdpx9b_inst_22_dout;
wire [26:0] sdpx9b_inst_23_dout_w;
wire [8:0] sdpx9b_inst_23_dout;
wire [26:0] sdpx9b_inst_24_dout_w;
wire [8:0] sdpx9b_inst_24_dout;
wire [26:0] sdpx9b_inst_25_dout_w;
wire [8:0] sdpx9b_inst_25_dout;
wire [26:0] sdpx9b_inst_26_dout_w;
wire [8:0] sdpx9b_inst_26_dout;
wire [26:0] sdpx9b_inst_27_dout_w;
wire [8:0] sdpx9b_inst_27_dout;
wire [26:0] sdpx9b_inst_28_dout_w;
wire [8:0] sdpx9b_inst_28_dout;
wire [26:0] sdpx9b_inst_29_dout_w;
wire [8:0] sdpx9b_inst_29_dout;
wire [26:0] sdpx9b_inst_30_dout_w;
wire [8:0] sdpx9b_inst_30_dout;
wire [26:0] sdpx9b_inst_31_dout_w;
wire [8:0] sdpx9b_inst_31_dout;
wire [30:0] sdpb_inst_32_dout_w;
wire [9:9] sdpb_inst_32_dout;
wire [30:0] sdpb_inst_33_dout_w;
wire [9:9] sdpb_inst_33_dout;
wire [30:0] sdpb_inst_34_dout_w;
wire [9:9] sdpb_inst_34_dout;
wire [30:0] sdpb_inst_35_dout_w;
wire [9:9] sdpb_inst_35_dout;
wire [30:0] sdpb_inst_36_dout_w;
wire [10:10] sdpb_inst_36_dout;
wire [30:0] sdpb_inst_37_dout_w;
wire [10:10] sdpb_inst_37_dout;
wire [30:0] sdpb_inst_38_dout_w;
wire [10:10] sdpb_inst_38_dout;
wire [30:0] sdpb_inst_39_dout_w;
wire [10:10] sdpb_inst_39_dout;
wire [30:0] sdpb_inst_40_dout_w;
wire [11:11] sdpb_inst_40_dout;
wire [30:0] sdpb_inst_41_dout_w;
wire [11:11] sdpb_inst_41_dout;
wire [30:0] sdpb_inst_42_dout_w;
wire [11:11] sdpb_inst_42_dout;
wire [30:0] sdpb_inst_43_dout_w;
wire [11:11] sdpb_inst_43_dout;
wire [30:0] sdpb_inst_44_dout_w;
wire [12:12] sdpb_inst_44_dout;
wire [30:0] sdpb_inst_45_dout_w;
wire [12:12] sdpb_inst_45_dout;
wire [30:0] sdpb_inst_46_dout_w;
wire [12:12] sdpb_inst_46_dout;
wire [30:0] sdpb_inst_47_dout_w;
wire [12:12] sdpb_inst_47_dout;
wire [30:0] sdpb_inst_48_dout_w;
wire [13:13] sdpb_inst_48_dout;
wire [30:0] sdpb_inst_49_dout_w;
wire [13:13] sdpb_inst_49_dout;
wire [30:0] sdpb_inst_50_dout_w;
wire [13:13] sdpb_inst_50_dout;
wire [30:0] sdpb_inst_51_dout_w;
wire [13:13] sdpb_inst_51_dout;
wire [30:0] sdpb_inst_52_dout_w;
wire [14:14] sdpb_inst_52_dout;
wire [30:0] sdpb_inst_53_dout_w;
wire [14:14] sdpb_inst_53_dout;
wire [30:0] sdpb_inst_54_dout_w;
wire [14:14] sdpb_inst_54_dout;
wire [30:0] sdpb_inst_55_dout_w;
wire [14:14] sdpb_inst_55_dout;
wire [30:0] sdpb_inst_56_dout_w;
wire [15:15] sdpb_inst_56_dout;
wire [30:0] sdpb_inst_57_dout_w;
wire [15:15] sdpb_inst_57_dout;
wire [30:0] sdpb_inst_58_dout_w;
wire [15:15] sdpb_inst_58_dout;
wire [30:0] sdpb_inst_59_dout_w;
wire [15:15] sdpb_inst_59_dout;
wire [26:0] sdpx9b_inst_60_dout_w;
wire [8:0] sdpx9b_inst_60_dout;
wire [26:0] sdpx9b_inst_61_dout_w;
wire [8:0] sdpx9b_inst_61_dout;
wire [26:0] sdpx9b_inst_62_dout_w;
wire [8:0] sdpx9b_inst_62_dout;
wire [26:0] sdpx9b_inst_63_dout_w;
wire [8:0] sdpx9b_inst_63_dout;
wire [26:0] sdpx9b_inst_64_dout_w;
wire [8:0] sdpx9b_inst_64_dout;
wire [26:0] sdpx9b_inst_65_dout_w;
wire [8:0] sdpx9b_inst_65_dout;
wire [26:0] sdpx9b_inst_66_dout_w;
wire [8:0] sdpx9b_inst_66_dout;
wire [26:0] sdpx9b_inst_67_dout_w;
wire [8:0] sdpx9b_inst_67_dout;
wire [26:0] sdpx9b_inst_68_dout_w;
wire [8:0] sdpx9b_inst_68_dout;
wire [26:0] sdpx9b_inst_69_dout_w;
wire [8:0] sdpx9b_inst_69_dout;
wire [26:0] sdpx9b_inst_70_dout_w;
wire [8:0] sdpx9b_inst_70_dout;
wire [26:0] sdpx9b_inst_71_dout_w;
wire [8:0] sdpx9b_inst_71_dout;
wire [26:0] sdpx9b_inst_72_dout_w;
wire [8:0] sdpx9b_inst_72_dout;
wire [26:0] sdpx9b_inst_73_dout_w;
wire [8:0] sdpx9b_inst_73_dout;
wire [26:0] sdpx9b_inst_74_dout_w;
wire [8:0] sdpx9b_inst_74_dout;
wire [26:0] sdpx9b_inst_75_dout_w;
wire [8:0] sdpx9b_inst_75_dout;
wire [30:0] sdpb_inst_76_dout_w;
wire [9:9] sdpb_inst_76_dout;
wire [30:0] sdpb_inst_77_dout_w;
wire [9:9] sdpb_inst_77_dout;
wire [30:0] sdpb_inst_78_dout_w;
wire [10:10] sdpb_inst_78_dout;
wire [30:0] sdpb_inst_79_dout_w;
wire [10:10] sdpb_inst_79_dout;
wire [30:0] sdpb_inst_80_dout_w;
wire [11:11] sdpb_inst_80_dout;
wire [30:0] sdpb_inst_81_dout_w;
wire [11:11] sdpb_inst_81_dout;
wire [30:0] sdpb_inst_82_dout_w;
wire [12:12] sdpb_inst_82_dout;
wire [30:0] sdpb_inst_83_dout_w;
wire [12:12] sdpb_inst_83_dout;
wire [30:0] sdpb_inst_84_dout_w;
wire [13:13] sdpb_inst_84_dout;
wire [30:0] sdpb_inst_85_dout_w;
wire [13:13] sdpb_inst_85_dout;
wire [30:0] sdpb_inst_86_dout_w;
wire [14:14] sdpb_inst_86_dout;
wire [30:0] sdpb_inst_87_dout_w;
wire [14:14] sdpb_inst_87_dout;
wire [30:0] sdpb_inst_88_dout_w;
wire [15:15] sdpb_inst_88_dout;
wire [30:0] sdpb_inst_89_dout_w;
wire [15:15] sdpb_inst_89_dout;
wire [26:0] sdpx9b_inst_90_dout_w;
wire [8:0] sdpx9b_inst_90_dout;
wire [26:0] sdpx9b_inst_91_dout_w;
wire [8:0] sdpx9b_inst_91_dout;
wire [26:0] sdpx9b_inst_92_dout_w;
wire [8:0] sdpx9b_inst_92_dout;
wire [26:0] sdpx9b_inst_93_dout_w;
wire [8:0] sdpx9b_inst_93_dout;
wire [26:0] sdpx9b_inst_94_dout_w;
wire [8:0] sdpx9b_inst_94_dout;
wire [26:0] sdpx9b_inst_95_dout_w;
wire [8:0] sdpx9b_inst_95_dout;
wire [26:0] sdpx9b_inst_96_dout_w;
wire [8:0] sdpx9b_inst_96_dout;
wire [26:0] sdpx9b_inst_97_dout_w;
wire [8:0] sdpx9b_inst_97_dout;
wire [30:0] sdpb_inst_98_dout_w;
wire [9:9] sdpb_inst_98_dout;
wire [30:0] sdpb_inst_99_dout_w;
wire [10:10] sdpb_inst_99_dout;
wire [30:0] sdpb_inst_100_dout_w;
wire [11:11] sdpb_inst_100_dout;
wire [30:0] sdpb_inst_101_dout_w;
wire [12:12] sdpb_inst_101_dout;
wire [30:0] sdpb_inst_102_dout_w;
wire [13:13] sdpb_inst_102_dout;
wire [30:0] sdpb_inst_103_dout_w;
wire [14:14] sdpb_inst_103_dout;
wire [30:0] sdpb_inst_104_dout_w;
wire [15:15] sdpb_inst_104_dout;
wire [29:0] sdpb_inst_105_dout_w;
wire [1:0] sdpb_inst_105_dout;
wire [29:0] sdpb_inst_106_dout_w;
wire [3:2] sdpb_inst_106_dout;
wire [29:0] sdpb_inst_107_dout_w;
wire [5:4] sdpb_inst_107_dout;
wire [29:0] sdpb_inst_108_dout_w;
wire [7:6] sdpb_inst_108_dout;
wire [29:0] sdpb_inst_109_dout_w;
wire [9:8] sdpb_inst_109_dout;
wire [29:0] sdpb_inst_110_dout_w;
wire [11:10] sdpb_inst_110_dout;
wire [29:0] sdpb_inst_111_dout_w;
wire [13:12] sdpb_inst_111_dout;
wire [29:0] sdpb_inst_112_dout_w;
wire [15:14] sdpb_inst_112_dout;
wire [27:0] sdpb_inst_113_dout_w;
wire [3:0] sdpb_inst_113_dout;
wire [27:0] sdpb_inst_114_dout_w;
wire [7:4] sdpb_inst_114_dout;
wire [27:0] sdpb_inst_115_dout_w;
wire [11:8] sdpb_inst_115_dout;
wire [27:0] sdpb_inst_116_dout_w;
wire [15:12] sdpb_inst_116_dout;
wire [15:0] sdpb_inst_117_dout_w;
wire [15:0] sdpb_inst_117_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_347;
wire mux_o_348;
wire mux_o_349;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_356;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_426;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_433;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_440;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_453;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_460;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_464;
wire mux_o_465;
wire mux_o_466;
wire mux_o_468;
wire mux_o_469;
wire mux_o_470;
wire mux_o_471;
wire mux_o_472;
wire mux_o_473;
wire mux_o_474;
wire mux_o_475;
wire mux_o_476;
wire mux_o_477;
wire mux_o_478;
wire mux_o_479;
wire mux_o_480;
wire mux_o_481;
wire mux_o_482;
wire mux_o_543;
wire mux_o_544;
wire mux_o_545;
wire mux_o_546;
wire mux_o_547;
wire mux_o_548;
wire mux_o_549;
wire mux_o_550;
wire mux_o_551;
wire mux_o_552;
wire mux_o_553;
wire mux_o_554;
wire mux_o_555;
wire mux_o_556;
wire mux_o_557;
wire mux_o_558;
wire mux_o_559;
wire mux_o_560;
wire mux_o_561;
wire mux_o_562;
wire mux_o_563;
wire mux_o_564;
wire mux_o_565;
wire mux_o_566;
wire mux_o_567;
wire mux_o_568;
wire mux_o_569;
wire mux_o_570;
wire mux_o_574;
wire mux_o_575;
wire mux_o_576;
wire mux_o_577;
wire mux_o_578;
wire mux_o_579;
wire mux_o_580;
wire mux_o_581;
wire mux_o_582;
wire mux_o_583;
wire mux_o_584;
wire mux_o_585;
wire mux_o_586;
wire mux_o_587;
wire mux_o_589;
wire mux_o_590;
wire mux_o_591;
wire mux_o_592;
wire mux_o_593;
wire mux_o_594;
wire mux_o_595;
wire mux_o_596;
wire mux_o_597;
wire mux_o_598;
wire mux_o_599;
wire mux_o_600;
wire mux_o_601;
wire mux_o_602;
wire mux_o_603;
wire mux_o_664;
wire mux_o_665;
wire mux_o_666;
wire mux_o_667;
wire mux_o_668;
wire mux_o_669;
wire mux_o_670;
wire mux_o_671;
wire mux_o_672;
wire mux_o_673;
wire mux_o_674;
wire mux_o_675;
wire mux_o_676;
wire mux_o_677;
wire mux_o_678;
wire mux_o_679;
wire mux_o_680;
wire mux_o_681;
wire mux_o_682;
wire mux_o_683;
wire mux_o_684;
wire mux_o_685;
wire mux_o_686;
wire mux_o_687;
wire mux_o_688;
wire mux_o_689;
wire mux_o_690;
wire mux_o_691;
wire mux_o_695;
wire mux_o_696;
wire mux_o_697;
wire mux_o_698;
wire mux_o_699;
wire mux_o_700;
wire mux_o_701;
wire mux_o_702;
wire mux_o_703;
wire mux_o_704;
wire mux_o_705;
wire mux_o_706;
wire mux_o_707;
wire mux_o_708;
wire mux_o_710;
wire mux_o_711;
wire mux_o_712;
wire mux_o_713;
wire mux_o_714;
wire mux_o_715;
wire mux_o_716;
wire mux_o_717;
wire mux_o_718;
wire mux_o_719;
wire mux_o_720;
wire mux_o_721;
wire mux_o_722;
wire mux_o_723;
wire mux_o_724;
wire mux_o_785;
wire mux_o_786;
wire mux_o_787;
wire mux_o_788;
wire mux_o_789;
wire mux_o_790;
wire mux_o_791;
wire mux_o_792;
wire mux_o_793;
wire mux_o_794;
wire mux_o_795;
wire mux_o_796;
wire mux_o_797;
wire mux_o_798;
wire mux_o_799;
wire mux_o_800;
wire mux_o_801;
wire mux_o_802;
wire mux_o_803;
wire mux_o_804;
wire mux_o_805;
wire mux_o_806;
wire mux_o_807;
wire mux_o_808;
wire mux_o_809;
wire mux_o_810;
wire mux_o_811;
wire mux_o_812;
wire mux_o_816;
wire mux_o_817;
wire mux_o_818;
wire mux_o_819;
wire mux_o_820;
wire mux_o_821;
wire mux_o_822;
wire mux_o_823;
wire mux_o_824;
wire mux_o_825;
wire mux_o_826;
wire mux_o_827;
wire mux_o_828;
wire mux_o_829;
wire mux_o_831;
wire mux_o_832;
wire mux_o_833;
wire mux_o_834;
wire mux_o_835;
wire mux_o_836;
wire mux_o_837;
wire mux_o_838;
wire mux_o_839;
wire mux_o_840;
wire mux_o_841;
wire mux_o_842;
wire mux_o_843;
wire mux_o_844;
wire mux_o_845;
wire mux_o_906;
wire mux_o_907;
wire mux_o_908;
wire mux_o_909;
wire mux_o_910;
wire mux_o_911;
wire mux_o_912;
wire mux_o_913;
wire mux_o_914;
wire mux_o_915;
wire mux_o_916;
wire mux_o_917;
wire mux_o_918;
wire mux_o_919;
wire mux_o_920;
wire mux_o_921;
wire mux_o_922;
wire mux_o_923;
wire mux_o_924;
wire mux_o_925;
wire mux_o_926;
wire mux_o_927;
wire mux_o_928;
wire mux_o_929;
wire mux_o_930;
wire mux_o_931;
wire mux_o_932;
wire mux_o_933;
wire mux_o_937;
wire mux_o_938;
wire mux_o_939;
wire mux_o_940;
wire mux_o_941;
wire mux_o_942;
wire mux_o_943;
wire mux_o_944;
wire mux_o_945;
wire mux_o_946;
wire mux_o_947;
wire mux_o_948;
wire mux_o_949;
wire mux_o_950;
wire mux_o_952;
wire mux_o_953;
wire mux_o_954;
wire mux_o_955;
wire mux_o_956;
wire mux_o_957;
wire mux_o_958;
wire mux_o_959;
wire mux_o_960;
wire mux_o_961;
wire mux_o_962;
wire mux_o_963;
wire mux_o_964;
wire mux_o_965;
wire mux_o_966;
wire mux_o_1027;
wire mux_o_1028;
wire mux_o_1029;
wire mux_o_1030;
wire mux_o_1031;
wire mux_o_1032;
wire mux_o_1033;
wire mux_o_1034;
wire mux_o_1035;
wire mux_o_1036;
wire mux_o_1037;
wire mux_o_1038;
wire mux_o_1039;
wire mux_o_1040;
wire mux_o_1041;
wire mux_o_1042;
wire mux_o_1043;
wire mux_o_1044;
wire mux_o_1045;
wire mux_o_1046;
wire mux_o_1047;
wire mux_o_1048;
wire mux_o_1049;
wire mux_o_1050;
wire mux_o_1051;
wire mux_o_1052;
wire mux_o_1053;
wire mux_o_1054;
wire mux_o_1058;
wire mux_o_1059;
wire mux_o_1060;
wire mux_o_1061;
wire mux_o_1062;
wire mux_o_1063;
wire mux_o_1064;
wire mux_o_1065;
wire mux_o_1066;
wire mux_o_1067;
wire mux_o_1068;
wire mux_o_1069;
wire mux_o_1070;
wire mux_o_1071;
wire mux_o_1073;
wire mux_o_1074;
wire mux_o_1075;
wire mux_o_1076;
wire mux_o_1077;
wire mux_o_1078;
wire mux_o_1079;
wire mux_o_1080;
wire mux_o_1081;
wire mux_o_1082;
wire mux_o_1083;
wire mux_o_1084;
wire mux_o_1085;
wire mux_o_1086;
wire mux_o_1087;
wire mux_o_1117;
wire mux_o_1125;
wire mux_o_1126;
wire mux_o_1127;
wire mux_o_1128;
wire mux_o_1129;
wire mux_o_1130;
wire mux_o_1131;
wire mux_o_1161;
wire mux_o_1169;
wire mux_o_1170;
wire mux_o_1171;
wire mux_o_1172;
wire mux_o_1173;
wire mux_o_1174;
wire mux_o_1175;
wire mux_o_1205;
wire mux_o_1213;
wire mux_o_1214;
wire mux_o_1215;
wire mux_o_1216;
wire mux_o_1217;
wire mux_o_1218;
wire mux_o_1219;
wire mux_o_1249;
wire mux_o_1257;
wire mux_o_1258;
wire mux_o_1259;
wire mux_o_1260;
wire mux_o_1261;
wire mux_o_1262;
wire mux_o_1263;
wire mux_o_1293;
wire mux_o_1301;
wire mux_o_1302;
wire mux_o_1303;
wire mux_o_1304;
wire mux_o_1305;
wire mux_o_1306;
wire mux_o_1307;
wire mux_o_1337;
wire mux_o_1345;
wire mux_o_1346;
wire mux_o_1347;
wire mux_o_1348;
wire mux_o_1349;
wire mux_o_1350;
wire mux_o_1351;
wire mux_o_1381;
wire mux_o_1389;
wire mux_o_1390;
wire mux_o_1391;
wire mux_o_1392;
wire mux_o_1393;
wire mux_o_1394;
wire mux_o_1395;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

LUT6 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_0.INIT = 64'h0000000000000001;
LUT6 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_1.INIT = 64'h0000000000000002;
LUT6 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_2.INIT = 64'h0000000000000004;
LUT6 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_3.INIT = 64'h0000000000000008;
LUT6 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_4.INIT = 64'h0000000000000010;
LUT6 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_5.INIT = 64'h0000000000000020;
LUT6 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_6.INIT = 64'h0000000000000040;
LUT6 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_7.INIT = 64'h0000000000000080;
LUT6 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_8.INIT = 64'h0000000000000100;
LUT6 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_9.INIT = 64'h0000000000000200;
LUT6 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_10.INIT = 64'h0000000000000400;
LUT6 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_11.INIT = 64'h0000000000000800;
LUT6 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_12.INIT = 64'h0000000000001000;
LUT6 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_13.INIT = 64'h0000000000002000;
LUT6 lut_inst_14 (
  .F(lut_f_14),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_14.INIT = 64'h0000000000004000;
LUT6 lut_inst_15 (
  .F(lut_f_15),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_15.INIT = 64'h0000000000008000;
LUT6 lut_inst_16 (
  .F(lut_f_16),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_16.INIT = 64'h0000000000010000;
LUT6 lut_inst_17 (
  .F(lut_f_17),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_17.INIT = 64'h0000000000020000;
LUT6 lut_inst_18 (
  .F(lut_f_18),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_18.INIT = 64'h0000000000040000;
LUT6 lut_inst_19 (
  .F(lut_f_19),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_19.INIT = 64'h0000000000080000;
LUT6 lut_inst_20 (
  .F(lut_f_20),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_20.INIT = 64'h0000000000100000;
LUT6 lut_inst_21 (
  .F(lut_f_21),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_21.INIT = 64'h0000000000200000;
LUT6 lut_inst_22 (
  .F(lut_f_22),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_22.INIT = 64'h0000000000400000;
LUT6 lut_inst_23 (
  .F(lut_f_23),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_23.INIT = 64'h0000000000800000;
LUT6 lut_inst_24 (
  .F(lut_f_24),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_24.INIT = 64'h0000000001000000;
LUT6 lut_inst_25 (
  .F(lut_f_25),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_25.INIT = 64'h0000000002000000;
LUT6 lut_inst_26 (
  .F(lut_f_26),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_26.INIT = 64'h0000000004000000;
LUT6 lut_inst_27 (
  .F(lut_f_27),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_27.INIT = 64'h0000000008000000;
LUT6 lut_inst_28 (
  .F(lut_f_28),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_28.INIT = 64'h0000000010000000;
LUT6 lut_inst_29 (
  .F(lut_f_29),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_29.INIT = 64'h0000000020000000;
LUT6 lut_inst_30 (
  .F(lut_f_30),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_30.INIT = 64'h0000000040000000;
LUT6 lut_inst_31 (
  .F(lut_f_31),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_31.INIT = 64'h0000000080000000;
LUT6 lut_inst_32 (
  .F(lut_f_32),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_32.INIT = 64'h0000000100000000;
LUT6 lut_inst_33 (
  .F(lut_f_33),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_33.INIT = 64'h0000000200000000;
LUT6 lut_inst_34 (
  .F(lut_f_34),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_34.INIT = 64'h0000000400000000;
LUT6 lut_inst_35 (
  .F(lut_f_35),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_35.INIT = 64'h0000000800000000;
LUT6 lut_inst_36 (
  .F(lut_f_36),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_36.INIT = 64'h0000001000000000;
LUT6 lut_inst_37 (
  .F(lut_f_37),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_37.INIT = 64'h0000002000000000;
LUT6 lut_inst_38 (
  .F(lut_f_38),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_38.INIT = 64'h0000004000000000;
LUT6 lut_inst_39 (
  .F(lut_f_39),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_39.INIT = 64'h0000008000000000;
LUT6 lut_inst_40 (
  .F(lut_f_40),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_40.INIT = 64'h0000010000000000;
LUT6 lut_inst_41 (
  .F(lut_f_41),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_41.INIT = 64'h0000020000000000;
LUT6 lut_inst_42 (
  .F(lut_f_42),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_42.INIT = 64'h0000040000000000;
LUT6 lut_inst_43 (
  .F(lut_f_43),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_43.INIT = 64'h0000080000000000;
LUT6 lut_inst_44 (
  .F(lut_f_44),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_44.INIT = 64'h0000100000000000;
LUT6 lut_inst_45 (
  .F(lut_f_45),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_45.INIT = 64'h0000200000000000;
LUT6 lut_inst_46 (
  .F(lut_f_46),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_46.INIT = 64'h0000400000000000;
LUT6 lut_inst_47 (
  .F(lut_f_47),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_47.INIT = 64'h0000800000000000;
LUT6 lut_inst_48 (
  .F(lut_f_48),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_48.INIT = 64'h0001000000000000;
LUT6 lut_inst_49 (
  .F(lut_f_49),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_49.INIT = 64'h0002000000000000;
LUT6 lut_inst_50 (
  .F(lut_f_50),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_50.INIT = 64'h0004000000000000;
LUT6 lut_inst_51 (
  .F(lut_f_51),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_51.INIT = 64'h0008000000000000;
LUT6 lut_inst_52 (
  .F(lut_f_52),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_52.INIT = 64'h0010000000000000;
LUT6 lut_inst_53 (
  .F(lut_f_53),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_53.INIT = 64'h0020000000000000;
LUT6 lut_inst_54 (
  .F(lut_f_54),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_54.INIT = 64'h0040000000000000;
LUT6 lut_inst_55 (
  .F(lut_f_55),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_55.INIT = 64'h0080000000000000;
LUT4 lut_inst_56 (
  .F(lut_f_56),
  .I0(ada[13]),
  .I1(ada[14]),
  .I2(ada[15]),
  .I3(ada[16])
);
defparam lut_inst_56.INIT = 16'h4000;
LUT5 lut_inst_57 (
  .F(lut_f_57),
  .I0(ada[12]),
  .I1(ada[13]),
  .I2(ada[14]),
  .I3(ada[15]),
  .I4(ada[16])
);
defparam lut_inst_57.INIT = 32'h40000000;
LUT7 lut_inst_58 (
  .F(lut_f_58),
  .I0(ada[10]),
  .I1(ada[11]),
  .I2(ada[12]),
  .I3(ada[13]),
  .I4(ada[14]),
  .I5(ada[15]),
  .I6(ada[16])
);
defparam lut_inst_58.INIT = 128'h10000000000000000000000000000000;
LUT6 lut_inst_59 (
  .F(lut_f_59),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_59.INIT = 64'h0000000000000001;
LUT6 lut_inst_60 (
  .F(lut_f_60),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_60.INIT = 64'h0000000000000002;
LUT6 lut_inst_61 (
  .F(lut_f_61),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_61.INIT = 64'h0000000000000004;
LUT6 lut_inst_62 (
  .F(lut_f_62),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_62.INIT = 64'h0000000000000008;
LUT6 lut_inst_63 (
  .F(lut_f_63),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_63.INIT = 64'h0000000000000010;
LUT6 lut_inst_64 (
  .F(lut_f_64),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_64.INIT = 64'h0000000000000020;
LUT6 lut_inst_65 (
  .F(lut_f_65),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_65.INIT = 64'h0000000000000040;
LUT6 lut_inst_66 (
  .F(lut_f_66),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_66.INIT = 64'h0000000000000080;
LUT6 lut_inst_67 (
  .F(lut_f_67),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_67.INIT = 64'h0000000000000100;
LUT6 lut_inst_68 (
  .F(lut_f_68),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_68.INIT = 64'h0000000000000200;
LUT6 lut_inst_69 (
  .F(lut_f_69),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_69.INIT = 64'h0000000000000400;
LUT6 lut_inst_70 (
  .F(lut_f_70),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_70.INIT = 64'h0000000000000800;
LUT6 lut_inst_71 (
  .F(lut_f_71),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_71.INIT = 64'h0000000000001000;
LUT6 lut_inst_72 (
  .F(lut_f_72),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_72.INIT = 64'h0000000000002000;
LUT6 lut_inst_73 (
  .F(lut_f_73),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_73.INIT = 64'h0000000000004000;
LUT6 lut_inst_74 (
  .F(lut_f_74),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_74.INIT = 64'h0000000000008000;
LUT6 lut_inst_75 (
  .F(lut_f_75),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_75.INIT = 64'h0000000000010000;
LUT6 lut_inst_76 (
  .F(lut_f_76),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_76.INIT = 64'h0000000000020000;
LUT6 lut_inst_77 (
  .F(lut_f_77),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_77.INIT = 64'h0000000000040000;
LUT6 lut_inst_78 (
  .F(lut_f_78),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_78.INIT = 64'h0000000000080000;
LUT6 lut_inst_79 (
  .F(lut_f_79),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_79.INIT = 64'h0000000000100000;
LUT6 lut_inst_80 (
  .F(lut_f_80),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_80.INIT = 64'h0000000000200000;
LUT6 lut_inst_81 (
  .F(lut_f_81),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_81.INIT = 64'h0000000000400000;
LUT6 lut_inst_82 (
  .F(lut_f_82),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_82.INIT = 64'h0000000000800000;
LUT6 lut_inst_83 (
  .F(lut_f_83),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_83.INIT = 64'h0000000001000000;
LUT6 lut_inst_84 (
  .F(lut_f_84),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_84.INIT = 64'h0000000002000000;
LUT6 lut_inst_85 (
  .F(lut_f_85),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_85.INIT = 64'h0000000004000000;
LUT6 lut_inst_86 (
  .F(lut_f_86),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_86.INIT = 64'h0000000008000000;
LUT6 lut_inst_87 (
  .F(lut_f_87),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_87.INIT = 64'h0000000010000000;
LUT6 lut_inst_88 (
  .F(lut_f_88),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_88.INIT = 64'h0000000020000000;
LUT6 lut_inst_89 (
  .F(lut_f_89),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_89.INIT = 64'h0000000040000000;
LUT6 lut_inst_90 (
  .F(lut_f_90),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_90.INIT = 64'h0000000080000000;
LUT6 lut_inst_91 (
  .F(lut_f_91),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_91.INIT = 64'h0000000100000000;
LUT6 lut_inst_92 (
  .F(lut_f_92),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_92.INIT = 64'h0000000200000000;
LUT6 lut_inst_93 (
  .F(lut_f_93),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_93.INIT = 64'h0000000400000000;
LUT6 lut_inst_94 (
  .F(lut_f_94),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_94.INIT = 64'h0000000800000000;
LUT6 lut_inst_95 (
  .F(lut_f_95),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_95.INIT = 64'h0000001000000000;
LUT6 lut_inst_96 (
  .F(lut_f_96),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_96.INIT = 64'h0000002000000000;
LUT6 lut_inst_97 (
  .F(lut_f_97),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_97.INIT = 64'h0000004000000000;
LUT6 lut_inst_98 (
  .F(lut_f_98),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_98.INIT = 64'h0000008000000000;
LUT6 lut_inst_99 (
  .F(lut_f_99),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_99.INIT = 64'h0000010000000000;
LUT6 lut_inst_100 (
  .F(lut_f_100),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_100.INIT = 64'h0000020000000000;
LUT6 lut_inst_101 (
  .F(lut_f_101),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_101.INIT = 64'h0000040000000000;
LUT6 lut_inst_102 (
  .F(lut_f_102),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_102.INIT = 64'h0000080000000000;
LUT6 lut_inst_103 (
  .F(lut_f_103),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_103.INIT = 64'h0000100000000000;
LUT6 lut_inst_104 (
  .F(lut_f_104),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_104.INIT = 64'h0000200000000000;
LUT6 lut_inst_105 (
  .F(lut_f_105),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_105.INIT = 64'h0000400000000000;
LUT6 lut_inst_106 (
  .F(lut_f_106),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_106.INIT = 64'h0000800000000000;
LUT6 lut_inst_107 (
  .F(lut_f_107),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_107.INIT = 64'h0001000000000000;
LUT6 lut_inst_108 (
  .F(lut_f_108),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_108.INIT = 64'h0002000000000000;
LUT6 lut_inst_109 (
  .F(lut_f_109),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_109.INIT = 64'h0004000000000000;
LUT6 lut_inst_110 (
  .F(lut_f_110),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_110.INIT = 64'h0008000000000000;
LUT6 lut_inst_111 (
  .F(lut_f_111),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_111.INIT = 64'h0010000000000000;
LUT6 lut_inst_112 (
  .F(lut_f_112),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_112.INIT = 64'h0020000000000000;
LUT6 lut_inst_113 (
  .F(lut_f_113),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_113.INIT = 64'h0040000000000000;
LUT6 lut_inst_114 (
  .F(lut_f_114),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_114.INIT = 64'h0080000000000000;
LUT4 lut_inst_115 (
  .F(lut_f_115),
  .I0(adb[13]),
  .I1(adb[14]),
  .I2(adb[15]),
  .I3(adb[16])
);
defparam lut_inst_115.INIT = 16'h4000;
LUT5 lut_inst_116 (
  .F(lut_f_116),
  .I0(adb[12]),
  .I1(adb[13]),
  .I2(adb[14]),
  .I3(adb[15]),
  .I4(adb[16])
);
defparam lut_inst_116.INIT = 32'h40000000;
LUT7 lut_inst_117 (
  .F(lut_f_117),
  .I0(adb[10]),
  .I1(adb[11]),
  .I2(adb[12]),
  .I3(adb[13]),
  .I4(adb[14]),
  .I5(adb[15]),
  .I6(adb[16])
);
defparam lut_inst_117.INIT = 128'h10000000000000000000000000000000;
SDPX9B sdpx9b_inst_0 (
    .DO({sdpx9b_inst_0_dout_w[26:0],sdpx9b_inst_0_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_59}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_0.READ_MODE = 1'b0;
defparam sdpx9b_inst_0.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_0.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_0.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_0.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_0.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_1 (
    .DO({sdpx9b_inst_1_dout_w[26:0],sdpx9b_inst_1_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_60}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_1.READ_MODE = 1'b0;
defparam sdpx9b_inst_1.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_1.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_1.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_2 (
    .DO({sdpx9b_inst_2_dout_w[26:0],sdpx9b_inst_2_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_61}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_2.READ_MODE = 1'b0;
defparam sdpx9b_inst_2.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_2.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_2.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_2.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_2.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_3 (
    .DO({sdpx9b_inst_3_dout_w[26:0],sdpx9b_inst_3_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_62}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_3.READ_MODE = 1'b0;
defparam sdpx9b_inst_3.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_3.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_3.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_4 (
    .DO({sdpx9b_inst_4_dout_w[26:0],sdpx9b_inst_4_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_63}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_4.READ_MODE = 1'b0;
defparam sdpx9b_inst_4.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_4.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_4.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_4.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_4.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_5 (
    .DO({sdpx9b_inst_5_dout_w[26:0],sdpx9b_inst_5_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_64}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_5.READ_MODE = 1'b0;
defparam sdpx9b_inst_5.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_5.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_5.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_6 (
    .DO({sdpx9b_inst_6_dout_w[26:0],sdpx9b_inst_6_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_65}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_6.READ_MODE = 1'b0;
defparam sdpx9b_inst_6.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_6.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_6.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_7 (
    .DO({sdpx9b_inst_7_dout_w[26:0],sdpx9b_inst_7_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_66}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_7.READ_MODE = 1'b0;
defparam sdpx9b_inst_7.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_7.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_7.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_8 (
    .DO({sdpx9b_inst_8_dout_w[26:0],sdpx9b_inst_8_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_67}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_8.READ_MODE = 1'b0;
defparam sdpx9b_inst_8.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_8.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_8.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_9 (
    .DO({sdpx9b_inst_9_dout_w[26:0],sdpx9b_inst_9_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_68}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_9.READ_MODE = 1'b0;
defparam sdpx9b_inst_9.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_9.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_9.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_10 (
    .DO({sdpx9b_inst_10_dout_w[26:0],sdpx9b_inst_10_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_69}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_10.READ_MODE = 1'b0;
defparam sdpx9b_inst_10.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_10.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_10.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_10.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_10.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_11 (
    .DO({sdpx9b_inst_11_dout_w[26:0],sdpx9b_inst_11_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_70}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_11.READ_MODE = 1'b0;
defparam sdpx9b_inst_11.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_11.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_11.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_11.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_11.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_12 (
    .DO({sdpx9b_inst_12_dout_w[26:0],sdpx9b_inst_12_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_71}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_12.READ_MODE = 1'b0;
defparam sdpx9b_inst_12.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_12.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_12.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_12.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_12.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_13 (
    .DO({sdpx9b_inst_13_dout_w[26:0],sdpx9b_inst_13_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_72}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_13.READ_MODE = 1'b0;
defparam sdpx9b_inst_13.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_13.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_13.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_14 (
    .DO({sdpx9b_inst_14_dout_w[26:0],sdpx9b_inst_14_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_73}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_14.READ_MODE = 1'b0;
defparam sdpx9b_inst_14.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_14.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_14.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_15 (
    .DO({sdpx9b_inst_15_dout_w[26:0],sdpx9b_inst_15_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_15}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_74}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_15.READ_MODE = 1'b0;
defparam sdpx9b_inst_15.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_15.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_15.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_15.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_15.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_16 (
    .DO({sdpx9b_inst_16_dout_w[26:0],sdpx9b_inst_16_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_16}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_75}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_16.READ_MODE = 1'b0;
defparam sdpx9b_inst_16.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_16.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_16.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_16.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_16.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_17 (
    .DO({sdpx9b_inst_17_dout_w[26:0],sdpx9b_inst_17_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_17}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_76}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_17.READ_MODE = 1'b0;
defparam sdpx9b_inst_17.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_17.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_17.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_17.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_17.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_18 (
    .DO({sdpx9b_inst_18_dout_w[26:0],sdpx9b_inst_18_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_18}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_77}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_18.READ_MODE = 1'b0;
defparam sdpx9b_inst_18.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_18.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_18.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_18.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_18.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_19 (
    .DO({sdpx9b_inst_19_dout_w[26:0],sdpx9b_inst_19_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_19}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_78}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_19.READ_MODE = 1'b0;
defparam sdpx9b_inst_19.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_19.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_19.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_19.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_19.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_20 (
    .DO({sdpx9b_inst_20_dout_w[26:0],sdpx9b_inst_20_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_20}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_79}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_20.READ_MODE = 1'b0;
defparam sdpx9b_inst_20.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_20.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_20.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_20.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_20.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_21 (
    .DO({sdpx9b_inst_21_dout_w[26:0],sdpx9b_inst_21_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_21}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_80}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_21.READ_MODE = 1'b0;
defparam sdpx9b_inst_21.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_21.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_21.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_21.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_21.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_22 (
    .DO({sdpx9b_inst_22_dout_w[26:0],sdpx9b_inst_22_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_22}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_81}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_22.READ_MODE = 1'b0;
defparam sdpx9b_inst_22.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_22.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_22.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_22.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_22.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_23 (
    .DO({sdpx9b_inst_23_dout_w[26:0],sdpx9b_inst_23_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_23}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_82}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_23.READ_MODE = 1'b0;
defparam sdpx9b_inst_23.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_23.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_23.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_23.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_23.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_24 (
    .DO({sdpx9b_inst_24_dout_w[26:0],sdpx9b_inst_24_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_24}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_83}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_24.READ_MODE = 1'b0;
defparam sdpx9b_inst_24.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_24.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_24.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_24.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_24.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_25 (
    .DO({sdpx9b_inst_25_dout_w[26:0],sdpx9b_inst_25_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_25}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_84}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_25.READ_MODE = 1'b0;
defparam sdpx9b_inst_25.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_25.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_25.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_25.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_25.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_26 (
    .DO({sdpx9b_inst_26_dout_w[26:0],sdpx9b_inst_26_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_26}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_85}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_26.READ_MODE = 1'b0;
defparam sdpx9b_inst_26.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_26.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_26.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_26.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_26.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_27 (
    .DO({sdpx9b_inst_27_dout_w[26:0],sdpx9b_inst_27_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_27}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_86}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_27.READ_MODE = 1'b0;
defparam sdpx9b_inst_27.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_27.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_27.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_27.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_27.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_28 (
    .DO({sdpx9b_inst_28_dout_w[26:0],sdpx9b_inst_28_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_28}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_87}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_28.READ_MODE = 1'b0;
defparam sdpx9b_inst_28.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_28.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_28.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_28.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_28.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_29 (
    .DO({sdpx9b_inst_29_dout_w[26:0],sdpx9b_inst_29_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_29}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_88}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_29.READ_MODE = 1'b0;
defparam sdpx9b_inst_29.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_29.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_29.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_29.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_29.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_30 (
    .DO({sdpx9b_inst_30_dout_w[26:0],sdpx9b_inst_30_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_30}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_89}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_30.READ_MODE = 1'b0;
defparam sdpx9b_inst_30.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_30.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_30.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_30.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_30.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_31 (
    .DO({sdpx9b_inst_31_dout_w[26:0],sdpx9b_inst_31_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_31}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_90}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_31.READ_MODE = 1'b0;
defparam sdpx9b_inst_31.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_31.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_31.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_31.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_31.RESET_MODE = "SYNC";

SDPB sdpb_inst_32 (
    .DO({sdpb_inst_32_dout_w[30:0],sdpb_inst_32_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_32.READ_MODE = 1'b0;
defparam sdpb_inst_32.BIT_WIDTH_0 = 1;
defparam sdpb_inst_32.BIT_WIDTH_1 = 1;
defparam sdpb_inst_32.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_32.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_32.RESET_MODE = "SYNC";

SDPB sdpb_inst_33 (
    .DO({sdpb_inst_33_dout_w[30:0],sdpb_inst_33_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_33.READ_MODE = 1'b0;
defparam sdpb_inst_33.BIT_WIDTH_0 = 1;
defparam sdpb_inst_33.BIT_WIDTH_1 = 1;
defparam sdpb_inst_33.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_33.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_33.RESET_MODE = "SYNC";

SDPB sdpb_inst_34 (
    .DO({sdpb_inst_34_dout_w[30:0],sdpb_inst_34_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_34.READ_MODE = 1'b0;
defparam sdpb_inst_34.BIT_WIDTH_0 = 1;
defparam sdpb_inst_34.BIT_WIDTH_1 = 1;
defparam sdpb_inst_34.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_34.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_34.RESET_MODE = "SYNC";

SDPB sdpb_inst_35 (
    .DO({sdpb_inst_35_dout_w[30:0],sdpb_inst_35_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_35.READ_MODE = 1'b0;
defparam sdpb_inst_35.BIT_WIDTH_0 = 1;
defparam sdpb_inst_35.BIT_WIDTH_1 = 1;
defparam sdpb_inst_35.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_35.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_35.RESET_MODE = "SYNC";

SDPB sdpb_inst_36 (
    .DO({sdpb_inst_36_dout_w[30:0],sdpb_inst_36_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_36.READ_MODE = 1'b0;
defparam sdpb_inst_36.BIT_WIDTH_0 = 1;
defparam sdpb_inst_36.BIT_WIDTH_1 = 1;
defparam sdpb_inst_36.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_36.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_36.RESET_MODE = "SYNC";

SDPB sdpb_inst_37 (
    .DO({sdpb_inst_37_dout_w[30:0],sdpb_inst_37_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_37.READ_MODE = 1'b0;
defparam sdpb_inst_37.BIT_WIDTH_0 = 1;
defparam sdpb_inst_37.BIT_WIDTH_1 = 1;
defparam sdpb_inst_37.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_37.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_37.RESET_MODE = "SYNC";

SDPB sdpb_inst_38 (
    .DO({sdpb_inst_38_dout_w[30:0],sdpb_inst_38_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_38.READ_MODE = 1'b0;
defparam sdpb_inst_38.BIT_WIDTH_0 = 1;
defparam sdpb_inst_38.BIT_WIDTH_1 = 1;
defparam sdpb_inst_38.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_38.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_38.RESET_MODE = "SYNC";

SDPB sdpb_inst_39 (
    .DO({sdpb_inst_39_dout_w[30:0],sdpb_inst_39_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_39.READ_MODE = 1'b0;
defparam sdpb_inst_39.BIT_WIDTH_0 = 1;
defparam sdpb_inst_39.BIT_WIDTH_1 = 1;
defparam sdpb_inst_39.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_39.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_39.RESET_MODE = "SYNC";

SDPB sdpb_inst_40 (
    .DO({sdpb_inst_40_dout_w[30:0],sdpb_inst_40_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_40.READ_MODE = 1'b0;
defparam sdpb_inst_40.BIT_WIDTH_0 = 1;
defparam sdpb_inst_40.BIT_WIDTH_1 = 1;
defparam sdpb_inst_40.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_40.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_40.RESET_MODE = "SYNC";

SDPB sdpb_inst_41 (
    .DO({sdpb_inst_41_dout_w[30:0],sdpb_inst_41_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_41.READ_MODE = 1'b0;
defparam sdpb_inst_41.BIT_WIDTH_0 = 1;
defparam sdpb_inst_41.BIT_WIDTH_1 = 1;
defparam sdpb_inst_41.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_41.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_41.RESET_MODE = "SYNC";

SDPB sdpb_inst_42 (
    .DO({sdpb_inst_42_dout_w[30:0],sdpb_inst_42_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_42.READ_MODE = 1'b0;
defparam sdpb_inst_42.BIT_WIDTH_0 = 1;
defparam sdpb_inst_42.BIT_WIDTH_1 = 1;
defparam sdpb_inst_42.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_42.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_42.RESET_MODE = "SYNC";

SDPB sdpb_inst_43 (
    .DO({sdpb_inst_43_dout_w[30:0],sdpb_inst_43_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_43.READ_MODE = 1'b0;
defparam sdpb_inst_43.BIT_WIDTH_0 = 1;
defparam sdpb_inst_43.BIT_WIDTH_1 = 1;
defparam sdpb_inst_43.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_43.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_43.RESET_MODE = "SYNC";

SDPB sdpb_inst_44 (
    .DO({sdpb_inst_44_dout_w[30:0],sdpb_inst_44_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_44.READ_MODE = 1'b0;
defparam sdpb_inst_44.BIT_WIDTH_0 = 1;
defparam sdpb_inst_44.BIT_WIDTH_1 = 1;
defparam sdpb_inst_44.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_44.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_44.RESET_MODE = "SYNC";

SDPB sdpb_inst_45 (
    .DO({sdpb_inst_45_dout_w[30:0],sdpb_inst_45_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_45.READ_MODE = 1'b0;
defparam sdpb_inst_45.BIT_WIDTH_0 = 1;
defparam sdpb_inst_45.BIT_WIDTH_1 = 1;
defparam sdpb_inst_45.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_45.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_45.RESET_MODE = "SYNC";

SDPB sdpb_inst_46 (
    .DO({sdpb_inst_46_dout_w[30:0],sdpb_inst_46_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_46.READ_MODE = 1'b0;
defparam sdpb_inst_46.BIT_WIDTH_0 = 1;
defparam sdpb_inst_46.BIT_WIDTH_1 = 1;
defparam sdpb_inst_46.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_46.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_46.RESET_MODE = "SYNC";

SDPB sdpb_inst_47 (
    .DO({sdpb_inst_47_dout_w[30:0],sdpb_inst_47_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_47.READ_MODE = 1'b0;
defparam sdpb_inst_47.BIT_WIDTH_0 = 1;
defparam sdpb_inst_47.BIT_WIDTH_1 = 1;
defparam sdpb_inst_47.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_47.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_47.RESET_MODE = "SYNC";

SDPB sdpb_inst_48 (
    .DO({sdpb_inst_48_dout_w[30:0],sdpb_inst_48_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_48.READ_MODE = 1'b0;
defparam sdpb_inst_48.BIT_WIDTH_0 = 1;
defparam sdpb_inst_48.BIT_WIDTH_1 = 1;
defparam sdpb_inst_48.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_48.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_48.RESET_MODE = "SYNC";

SDPB sdpb_inst_49 (
    .DO({sdpb_inst_49_dout_w[30:0],sdpb_inst_49_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_49.READ_MODE = 1'b0;
defparam sdpb_inst_49.BIT_WIDTH_0 = 1;
defparam sdpb_inst_49.BIT_WIDTH_1 = 1;
defparam sdpb_inst_49.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_49.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_49.RESET_MODE = "SYNC";

SDPB sdpb_inst_50 (
    .DO({sdpb_inst_50_dout_w[30:0],sdpb_inst_50_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_50.READ_MODE = 1'b0;
defparam sdpb_inst_50.BIT_WIDTH_0 = 1;
defparam sdpb_inst_50.BIT_WIDTH_1 = 1;
defparam sdpb_inst_50.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_50.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_50.RESET_MODE = "SYNC";

SDPB sdpb_inst_51 (
    .DO({sdpb_inst_51_dout_w[30:0],sdpb_inst_51_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_51.READ_MODE = 1'b0;
defparam sdpb_inst_51.BIT_WIDTH_0 = 1;
defparam sdpb_inst_51.BIT_WIDTH_1 = 1;
defparam sdpb_inst_51.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_51.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_51.RESET_MODE = "SYNC";

SDPB sdpb_inst_52 (
    .DO({sdpb_inst_52_dout_w[30:0],sdpb_inst_52_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_52.READ_MODE = 1'b0;
defparam sdpb_inst_52.BIT_WIDTH_0 = 1;
defparam sdpb_inst_52.BIT_WIDTH_1 = 1;
defparam sdpb_inst_52.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_52.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_52.RESET_MODE = "SYNC";

SDPB sdpb_inst_53 (
    .DO({sdpb_inst_53_dout_w[30:0],sdpb_inst_53_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_53.READ_MODE = 1'b0;
defparam sdpb_inst_53.BIT_WIDTH_0 = 1;
defparam sdpb_inst_53.BIT_WIDTH_1 = 1;
defparam sdpb_inst_53.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_53.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_53.RESET_MODE = "SYNC";

SDPB sdpb_inst_54 (
    .DO({sdpb_inst_54_dout_w[30:0],sdpb_inst_54_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_54.READ_MODE = 1'b0;
defparam sdpb_inst_54.BIT_WIDTH_0 = 1;
defparam sdpb_inst_54.BIT_WIDTH_1 = 1;
defparam sdpb_inst_54.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_54.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_54.RESET_MODE = "SYNC";

SDPB sdpb_inst_55 (
    .DO({sdpb_inst_55_dout_w[30:0],sdpb_inst_55_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_55.READ_MODE = 1'b0;
defparam sdpb_inst_55.BIT_WIDTH_0 = 1;
defparam sdpb_inst_55.BIT_WIDTH_1 = 1;
defparam sdpb_inst_55.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_55.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_55.RESET_MODE = "SYNC";

SDPB sdpb_inst_56 (
    .DO({sdpb_inst_56_dout_w[30:0],sdpb_inst_56_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_56.READ_MODE = 1'b0;
defparam sdpb_inst_56.BIT_WIDTH_0 = 1;
defparam sdpb_inst_56.BIT_WIDTH_1 = 1;
defparam sdpb_inst_56.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_56.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_56.RESET_MODE = "SYNC";

SDPB sdpb_inst_57 (
    .DO({sdpb_inst_57_dout_w[30:0],sdpb_inst_57_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_57.READ_MODE = 1'b0;
defparam sdpb_inst_57.BIT_WIDTH_0 = 1;
defparam sdpb_inst_57.BIT_WIDTH_1 = 1;
defparam sdpb_inst_57.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_57.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_57.RESET_MODE = "SYNC";

SDPB sdpb_inst_58 (
    .DO({sdpb_inst_58_dout_w[30:0],sdpb_inst_58_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_58.READ_MODE = 1'b0;
defparam sdpb_inst_58.BIT_WIDTH_0 = 1;
defparam sdpb_inst_58.BIT_WIDTH_1 = 1;
defparam sdpb_inst_58.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_58.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_58.RESET_MODE = "SYNC";

SDPB sdpb_inst_59 (
    .DO({sdpb_inst_59_dout_w[30:0],sdpb_inst_59_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_59.READ_MODE = 1'b0;
defparam sdpb_inst_59.BIT_WIDTH_0 = 1;
defparam sdpb_inst_59.BIT_WIDTH_1 = 1;
defparam sdpb_inst_59.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_59.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_59.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_60 (
    .DO({sdpx9b_inst_60_dout_w[26:0],sdpx9b_inst_60_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_32}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_91}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_60.READ_MODE = 1'b0;
defparam sdpx9b_inst_60.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_60.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_60.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_60.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_60.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_61 (
    .DO({sdpx9b_inst_61_dout_w[26:0],sdpx9b_inst_61_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_33}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_92}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_61.READ_MODE = 1'b0;
defparam sdpx9b_inst_61.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_61.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_61.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_61.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_61.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_62 (
    .DO({sdpx9b_inst_62_dout_w[26:0],sdpx9b_inst_62_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_34}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_93}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_62.READ_MODE = 1'b0;
defparam sdpx9b_inst_62.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_62.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_62.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_62.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_62.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_63 (
    .DO({sdpx9b_inst_63_dout_w[26:0],sdpx9b_inst_63_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_35}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_94}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_63.READ_MODE = 1'b0;
defparam sdpx9b_inst_63.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_63.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_63.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_63.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_63.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_64 (
    .DO({sdpx9b_inst_64_dout_w[26:0],sdpx9b_inst_64_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_36}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_95}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_64.READ_MODE = 1'b0;
defparam sdpx9b_inst_64.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_64.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_64.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_64.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_64.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_65 (
    .DO({sdpx9b_inst_65_dout_w[26:0],sdpx9b_inst_65_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_37}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_96}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_65.READ_MODE = 1'b0;
defparam sdpx9b_inst_65.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_65.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_65.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_65.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_65.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_66 (
    .DO({sdpx9b_inst_66_dout_w[26:0],sdpx9b_inst_66_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_38}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_97}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_66.READ_MODE = 1'b0;
defparam sdpx9b_inst_66.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_66.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_66.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_66.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_66.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_67 (
    .DO({sdpx9b_inst_67_dout_w[26:0],sdpx9b_inst_67_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_39}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_98}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_67.READ_MODE = 1'b0;
defparam sdpx9b_inst_67.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_67.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_67.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_67.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_67.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_68 (
    .DO({sdpx9b_inst_68_dout_w[26:0],sdpx9b_inst_68_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_40}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_99}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_68.READ_MODE = 1'b0;
defparam sdpx9b_inst_68.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_68.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_68.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_68.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_68.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_69 (
    .DO({sdpx9b_inst_69_dout_w[26:0],sdpx9b_inst_69_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_41}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_100}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_69.READ_MODE = 1'b0;
defparam sdpx9b_inst_69.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_69.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_69.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_69.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_69.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_70 (
    .DO({sdpx9b_inst_70_dout_w[26:0],sdpx9b_inst_70_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_42}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_101}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_70.READ_MODE = 1'b0;
defparam sdpx9b_inst_70.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_70.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_70.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_70.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_70.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_71 (
    .DO({sdpx9b_inst_71_dout_w[26:0],sdpx9b_inst_71_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_43}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_102}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_71.READ_MODE = 1'b0;
defparam sdpx9b_inst_71.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_71.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_71.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_71.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_71.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_72 (
    .DO({sdpx9b_inst_72_dout_w[26:0],sdpx9b_inst_72_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_44}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_103}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_72.READ_MODE = 1'b0;
defparam sdpx9b_inst_72.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_72.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_72.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_72.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_72.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_73 (
    .DO({sdpx9b_inst_73_dout_w[26:0],sdpx9b_inst_73_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_45}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_104}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_73.READ_MODE = 1'b0;
defparam sdpx9b_inst_73.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_73.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_73.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_73.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_73.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_74 (
    .DO({sdpx9b_inst_74_dout_w[26:0],sdpx9b_inst_74_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_46}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_105}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_74.READ_MODE = 1'b0;
defparam sdpx9b_inst_74.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_74.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_74.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_74.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_74.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_75 (
    .DO({sdpx9b_inst_75_dout_w[26:0],sdpx9b_inst_75_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_47}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_106}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_75.READ_MODE = 1'b0;
defparam sdpx9b_inst_75.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_75.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_75.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_75.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_75.RESET_MODE = "SYNC";

SDPB sdpb_inst_76 (
    .DO({sdpb_inst_76_dout_w[30:0],sdpb_inst_76_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_76.READ_MODE = 1'b0;
defparam sdpb_inst_76.BIT_WIDTH_0 = 1;
defparam sdpb_inst_76.BIT_WIDTH_1 = 1;
defparam sdpb_inst_76.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_76.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_76.RESET_MODE = "SYNC";

SDPB sdpb_inst_77 (
    .DO({sdpb_inst_77_dout_w[30:0],sdpb_inst_77_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_77.READ_MODE = 1'b0;
defparam sdpb_inst_77.BIT_WIDTH_0 = 1;
defparam sdpb_inst_77.BIT_WIDTH_1 = 1;
defparam sdpb_inst_77.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_77.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_77.RESET_MODE = "SYNC";

SDPB sdpb_inst_78 (
    .DO({sdpb_inst_78_dout_w[30:0],sdpb_inst_78_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_78.READ_MODE = 1'b0;
defparam sdpb_inst_78.BIT_WIDTH_0 = 1;
defparam sdpb_inst_78.BIT_WIDTH_1 = 1;
defparam sdpb_inst_78.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_78.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_78.RESET_MODE = "SYNC";

SDPB sdpb_inst_79 (
    .DO({sdpb_inst_79_dout_w[30:0],sdpb_inst_79_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_79.READ_MODE = 1'b0;
defparam sdpb_inst_79.BIT_WIDTH_0 = 1;
defparam sdpb_inst_79.BIT_WIDTH_1 = 1;
defparam sdpb_inst_79.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_79.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_79.RESET_MODE = "SYNC";

SDPB sdpb_inst_80 (
    .DO({sdpb_inst_80_dout_w[30:0],sdpb_inst_80_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_80.READ_MODE = 1'b0;
defparam sdpb_inst_80.BIT_WIDTH_0 = 1;
defparam sdpb_inst_80.BIT_WIDTH_1 = 1;
defparam sdpb_inst_80.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_80.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_80.RESET_MODE = "SYNC";

SDPB sdpb_inst_81 (
    .DO({sdpb_inst_81_dout_w[30:0],sdpb_inst_81_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_81.READ_MODE = 1'b0;
defparam sdpb_inst_81.BIT_WIDTH_0 = 1;
defparam sdpb_inst_81.BIT_WIDTH_1 = 1;
defparam sdpb_inst_81.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_81.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_81.RESET_MODE = "SYNC";

SDPB sdpb_inst_82 (
    .DO({sdpb_inst_82_dout_w[30:0],sdpb_inst_82_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_82.READ_MODE = 1'b0;
defparam sdpb_inst_82.BIT_WIDTH_0 = 1;
defparam sdpb_inst_82.BIT_WIDTH_1 = 1;
defparam sdpb_inst_82.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_82.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_82.RESET_MODE = "SYNC";

SDPB sdpb_inst_83 (
    .DO({sdpb_inst_83_dout_w[30:0],sdpb_inst_83_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_83.READ_MODE = 1'b0;
defparam sdpb_inst_83.BIT_WIDTH_0 = 1;
defparam sdpb_inst_83.BIT_WIDTH_1 = 1;
defparam sdpb_inst_83.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_83.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_83.RESET_MODE = "SYNC";

SDPB sdpb_inst_84 (
    .DO({sdpb_inst_84_dout_w[30:0],sdpb_inst_84_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_84.READ_MODE = 1'b0;
defparam sdpb_inst_84.BIT_WIDTH_0 = 1;
defparam sdpb_inst_84.BIT_WIDTH_1 = 1;
defparam sdpb_inst_84.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_84.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_84.RESET_MODE = "SYNC";

SDPB sdpb_inst_85 (
    .DO({sdpb_inst_85_dout_w[30:0],sdpb_inst_85_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_85.READ_MODE = 1'b0;
defparam sdpb_inst_85.BIT_WIDTH_0 = 1;
defparam sdpb_inst_85.BIT_WIDTH_1 = 1;
defparam sdpb_inst_85.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_85.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_85.RESET_MODE = "SYNC";

SDPB sdpb_inst_86 (
    .DO({sdpb_inst_86_dout_w[30:0],sdpb_inst_86_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_86.READ_MODE = 1'b0;
defparam sdpb_inst_86.BIT_WIDTH_0 = 1;
defparam sdpb_inst_86.BIT_WIDTH_1 = 1;
defparam sdpb_inst_86.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_86.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_86.RESET_MODE = "SYNC";

SDPB sdpb_inst_87 (
    .DO({sdpb_inst_87_dout_w[30:0],sdpb_inst_87_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_87.READ_MODE = 1'b0;
defparam sdpb_inst_87.BIT_WIDTH_0 = 1;
defparam sdpb_inst_87.BIT_WIDTH_1 = 1;
defparam sdpb_inst_87.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_87.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_87.RESET_MODE = "SYNC";

SDPB sdpb_inst_88 (
    .DO({sdpb_inst_88_dout_w[30:0],sdpb_inst_88_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_88.READ_MODE = 1'b0;
defparam sdpb_inst_88.BIT_WIDTH_0 = 1;
defparam sdpb_inst_88.BIT_WIDTH_1 = 1;
defparam sdpb_inst_88.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_88.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_88.RESET_MODE = "SYNC";

SDPB sdpb_inst_89 (
    .DO({sdpb_inst_89_dout_w[30:0],sdpb_inst_89_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_89.READ_MODE = 1'b0;
defparam sdpb_inst_89.BIT_WIDTH_0 = 1;
defparam sdpb_inst_89.BIT_WIDTH_1 = 1;
defparam sdpb_inst_89.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_89.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_89.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_90 (
    .DO({sdpx9b_inst_90_dout_w[26:0],sdpx9b_inst_90_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_48}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_107}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_90.READ_MODE = 1'b0;
defparam sdpx9b_inst_90.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_90.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_90.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_90.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_90.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_91 (
    .DO({sdpx9b_inst_91_dout_w[26:0],sdpx9b_inst_91_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_49}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_108}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_91.READ_MODE = 1'b0;
defparam sdpx9b_inst_91.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_91.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_91.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_91.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_91.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_92 (
    .DO({sdpx9b_inst_92_dout_w[26:0],sdpx9b_inst_92_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_50}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_109}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_92.READ_MODE = 1'b0;
defparam sdpx9b_inst_92.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_92.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_92.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_92.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_92.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_93 (
    .DO({sdpx9b_inst_93_dout_w[26:0],sdpx9b_inst_93_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_51}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_110}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_93.READ_MODE = 1'b0;
defparam sdpx9b_inst_93.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_93.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_93.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_93.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_93.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_94 (
    .DO({sdpx9b_inst_94_dout_w[26:0],sdpx9b_inst_94_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_52}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_111}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_94.READ_MODE = 1'b0;
defparam sdpx9b_inst_94.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_94.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_94.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_94.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_94.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_95 (
    .DO({sdpx9b_inst_95_dout_w[26:0],sdpx9b_inst_95_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_53}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_112}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_95.READ_MODE = 1'b0;
defparam sdpx9b_inst_95.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_95.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_95.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_95.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_95.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_96 (
    .DO({sdpx9b_inst_96_dout_w[26:0],sdpx9b_inst_96_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_54}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_113}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_96.READ_MODE = 1'b0;
defparam sdpx9b_inst_96.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_96.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_96.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_96.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_96.RESET_MODE = "SYNC";

SDPX9B sdpx9b_inst_97 (
    .DO({sdpx9b_inst_97_dout_w[26:0],sdpx9b_inst_97_dout[8:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_55}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_114}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpx9b_inst_97.READ_MODE = 1'b0;
defparam sdpx9b_inst_97.BIT_WIDTH_0 = 9;
defparam sdpx9b_inst_97.BIT_WIDTH_1 = 9;
defparam sdpx9b_inst_97.BLK_SEL_0 = 3'b001;
defparam sdpx9b_inst_97.BLK_SEL_1 = 3'b001;
defparam sdpx9b_inst_97.RESET_MODE = "SYNC";

SDPB sdpb_inst_98 (
    .DO({sdpb_inst_98_dout_w[30:0],sdpb_inst_98_dout[9]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_98.READ_MODE = 1'b0;
defparam sdpb_inst_98.BIT_WIDTH_0 = 1;
defparam sdpb_inst_98.BIT_WIDTH_1 = 1;
defparam sdpb_inst_98.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_98.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_98.RESET_MODE = "SYNC";

SDPB sdpb_inst_99 (
    .DO({sdpb_inst_99_dout_w[30:0],sdpb_inst_99_dout[10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_99.READ_MODE = 1'b0;
defparam sdpb_inst_99.BIT_WIDTH_0 = 1;
defparam sdpb_inst_99.BIT_WIDTH_1 = 1;
defparam sdpb_inst_99.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_99.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_99.RESET_MODE = "SYNC";

SDPB sdpb_inst_100 (
    .DO({sdpb_inst_100_dout_w[30:0],sdpb_inst_100_dout[11]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_100.READ_MODE = 1'b0;
defparam sdpb_inst_100.BIT_WIDTH_0 = 1;
defparam sdpb_inst_100.BIT_WIDTH_1 = 1;
defparam sdpb_inst_100.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_100.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_100.RESET_MODE = "SYNC";

SDPB sdpb_inst_101 (
    .DO({sdpb_inst_101_dout_w[30:0],sdpb_inst_101_dout[12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_101.READ_MODE = 1'b0;
defparam sdpb_inst_101.BIT_WIDTH_0 = 1;
defparam sdpb_inst_101.BIT_WIDTH_1 = 1;
defparam sdpb_inst_101.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_101.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_101.RESET_MODE = "SYNC";

SDPB sdpb_inst_102 (
    .DO({sdpb_inst_102_dout_w[30:0],sdpb_inst_102_dout[13]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_102.READ_MODE = 1'b0;
defparam sdpb_inst_102.BIT_WIDTH_0 = 1;
defparam sdpb_inst_102.BIT_WIDTH_1 = 1;
defparam sdpb_inst_102.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_102.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_102.RESET_MODE = "SYNC";

SDPB sdpb_inst_103 (
    .DO({sdpb_inst_103_dout_w[30:0],sdpb_inst_103_dout[14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_103.READ_MODE = 1'b0;
defparam sdpb_inst_103.BIT_WIDTH_0 = 1;
defparam sdpb_inst_103.BIT_WIDTH_1 = 1;
defparam sdpb_inst_103.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_103.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_103.RESET_MODE = "SYNC";

SDPB sdpb_inst_104 (
    .DO({sdpb_inst_104_dout_w[30:0],sdpb_inst_104_dout[15]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_104.READ_MODE = 1'b0;
defparam sdpb_inst_104.BIT_WIDTH_0 = 1;
defparam sdpb_inst_104.BIT_WIDTH_1 = 1;
defparam sdpb_inst_104.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_104.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_104.RESET_MODE = "SYNC";

SDPB sdpb_inst_105 (
    .DO({sdpb_inst_105_dout_w[29:0],sdpb_inst_105_dout[1:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_105.READ_MODE = 1'b0;
defparam sdpb_inst_105.BIT_WIDTH_0 = 2;
defparam sdpb_inst_105.BIT_WIDTH_1 = 2;
defparam sdpb_inst_105.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_105.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_105.RESET_MODE = "SYNC";

SDPB sdpb_inst_106 (
    .DO({sdpb_inst_106_dout_w[29:0],sdpb_inst_106_dout[3:2]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_106.READ_MODE = 1'b0;
defparam sdpb_inst_106.BIT_WIDTH_0 = 2;
defparam sdpb_inst_106.BIT_WIDTH_1 = 2;
defparam sdpb_inst_106.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_106.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_106.RESET_MODE = "SYNC";

SDPB sdpb_inst_107 (
    .DO({sdpb_inst_107_dout_w[29:0],sdpb_inst_107_dout[5:4]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_107.READ_MODE = 1'b0;
defparam sdpb_inst_107.BIT_WIDTH_0 = 2;
defparam sdpb_inst_107.BIT_WIDTH_1 = 2;
defparam sdpb_inst_107.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_107.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_107.RESET_MODE = "SYNC";

SDPB sdpb_inst_108 (
    .DO({sdpb_inst_108_dout_w[29:0],sdpb_inst_108_dout[7:6]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_108.READ_MODE = 1'b0;
defparam sdpb_inst_108.BIT_WIDTH_0 = 2;
defparam sdpb_inst_108.BIT_WIDTH_1 = 2;
defparam sdpb_inst_108.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_108.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_108.RESET_MODE = "SYNC";

SDPB sdpb_inst_109 (
    .DO({sdpb_inst_109_dout_w[29:0],sdpb_inst_109_dout[9:8]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9:8]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_109.READ_MODE = 1'b0;
defparam sdpb_inst_109.BIT_WIDTH_0 = 2;
defparam sdpb_inst_109.BIT_WIDTH_1 = 2;
defparam sdpb_inst_109.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_109.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_109.RESET_MODE = "SYNC";

SDPB sdpb_inst_110 (
    .DO({sdpb_inst_110_dout_w[29:0],sdpb_inst_110_dout[11:10]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11:10]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_110.READ_MODE = 1'b0;
defparam sdpb_inst_110.BIT_WIDTH_0 = 2;
defparam sdpb_inst_110.BIT_WIDTH_1 = 2;
defparam sdpb_inst_110.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_110.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_110.RESET_MODE = "SYNC";

SDPB sdpb_inst_111 (
    .DO({sdpb_inst_111_dout_w[29:0],sdpb_inst_111_dout[13:12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13:12]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_111.READ_MODE = 1'b0;
defparam sdpb_inst_111.BIT_WIDTH_0 = 2;
defparam sdpb_inst_111.BIT_WIDTH_1 = 2;
defparam sdpb_inst_111.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_111.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_111.RESET_MODE = "SYNC";

SDPB sdpb_inst_112 (
    .DO({sdpb_inst_112_dout_w[29:0],sdpb_inst_112_dout[15:14]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_56}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_115}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:14]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_112.READ_MODE = 1'b0;
defparam sdpb_inst_112.BIT_WIDTH_0 = 2;
defparam sdpb_inst_112.BIT_WIDTH_1 = 2;
defparam sdpb_inst_112.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_112.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_112.RESET_MODE = "SYNC";

SDPB sdpb_inst_113 (
    .DO({sdpb_inst_113_dout_w[27:0],sdpb_inst_113_dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_116}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_113.READ_MODE = 1'b0;
defparam sdpb_inst_113.BIT_WIDTH_0 = 4;
defparam sdpb_inst_113.BIT_WIDTH_1 = 4;
defparam sdpb_inst_113.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_113.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_113.RESET_MODE = "SYNC";

SDPB sdpb_inst_114 (
    .DO({sdpb_inst_114_dout_w[27:0],sdpb_inst_114_dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_116}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_114.READ_MODE = 1'b0;
defparam sdpb_inst_114.BIT_WIDTH_0 = 4;
defparam sdpb_inst_114.BIT_WIDTH_1 = 4;
defparam sdpb_inst_114.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_114.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_114.RESET_MODE = "SYNC";

SDPB sdpb_inst_115 (
    .DO({sdpb_inst_115_dout_w[27:0],sdpb_inst_115_dout[11:8]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_116}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11:8]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_115.READ_MODE = 1'b0;
defparam sdpb_inst_115.BIT_WIDTH_0 = 4;
defparam sdpb_inst_115.BIT_WIDTH_1 = 4;
defparam sdpb_inst_115.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_115.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_115.RESET_MODE = "SYNC";

SDPB sdpb_inst_116 (
    .DO({sdpb_inst_116_dout_w[27:0],sdpb_inst_116_dout[15:12]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_57}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_116}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:12]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_116.READ_MODE = 1'b0;
defparam sdpb_inst_116.BIT_WIDTH_0 = 4;
defparam sdpb_inst_116.BIT_WIDTH_1 = 4;
defparam sdpb_inst_116.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_116.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_116.RESET_MODE = "SYNC";

SDPB sdpb_inst_117 (
    .DO({sdpb_inst_117_dout_w[15:0],sdpb_inst_117_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .CLKB(clkb),
    .CEB(ceb),
    .OCE(oce),
    .RESET(reset),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_58}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_117}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_117.READ_MODE = 1'b0;
defparam sdpb_inst_117.BIT_WIDTH_0 = 16;
defparam sdpb_inst_117.BIT_WIDTH_1 = 16;
defparam sdpb_inst_117.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_117.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_117.RESET_MODE = "SYNC";

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[16]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
DFFRE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb),
  .RESET(gw_gnd)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(sdpx9b_inst_0_dout[0]),
  .I1(sdpx9b_inst_1_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(sdpx9b_inst_2_dout[0]),
  .I1(sdpx9b_inst_3_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(sdpx9b_inst_4_dout[0]),
  .I1(sdpx9b_inst_5_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(sdpx9b_inst_6_dout[0]),
  .I1(sdpx9b_inst_7_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(sdpx9b_inst_8_dout[0]),
  .I1(sdpx9b_inst_9_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(sdpx9b_inst_10_dout[0]),
  .I1(sdpx9b_inst_11_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(sdpx9b_inst_12_dout[0]),
  .I1(sdpx9b_inst_13_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sdpx9b_inst_14_dout[0]),
  .I1(sdpx9b_inst_15_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sdpx9b_inst_16_dout[0]),
  .I1(sdpx9b_inst_17_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(sdpx9b_inst_18_dout[0]),
  .I1(sdpx9b_inst_19_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(sdpx9b_inst_20_dout[0]),
  .I1(sdpx9b_inst_21_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(sdpx9b_inst_22_dout[0]),
  .I1(sdpx9b_inst_23_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(sdpx9b_inst_24_dout[0]),
  .I1(sdpx9b_inst_25_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(sdpx9b_inst_26_dout[0]),
  .I1(sdpx9b_inst_27_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(sdpx9b_inst_28_dout[0]),
  .I1(sdpx9b_inst_29_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(sdpx9b_inst_30_dout[0]),
  .I1(sdpx9b_inst_31_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(sdpx9b_inst_60_dout[0]),
  .I1(sdpx9b_inst_61_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sdpx9b_inst_62_dout[0]),
  .I1(sdpx9b_inst_63_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(sdpx9b_inst_64_dout[0]),
  .I1(sdpx9b_inst_65_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sdpx9b_inst_66_dout[0]),
  .I1(sdpx9b_inst_67_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(sdpx9b_inst_68_dout[0]),
  .I1(sdpx9b_inst_69_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(sdpx9b_inst_70_dout[0]),
  .I1(sdpx9b_inst_71_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(sdpx9b_inst_72_dout[0]),
  .I1(sdpx9b_inst_73_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(sdpx9b_inst_74_dout[0]),
  .I1(sdpx9b_inst_75_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(sdpx9b_inst_90_dout[0]),
  .I1(sdpx9b_inst_91_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(sdpx9b_inst_92_dout[0]),
  .I1(sdpx9b_inst_93_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(sdpx9b_inst_94_dout[0]),
  .I1(sdpx9b_inst_95_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(sdpx9b_inst_96_dout[0]),
  .I1(sdpx9b_inst_97_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_59),
  .I1(mux_o_60),
  .S0(dff_q_4)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_61),
  .I1(mux_o_62),
  .S0(dff_q_4)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_63),
  .I1(mux_o_64),
  .S0(dff_q_4)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_65),
  .I1(mux_o_66),
  .S0(dff_q_4)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(mux_o_67),
  .I1(mux_o_68),
  .S0(dff_q_4)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_69),
  .I1(mux_o_70),
  .S0(dff_q_4)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_71),
  .I1(mux_o_72),
  .S0(dff_q_4)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_73),
  .I1(mux_o_74),
  .S0(dff_q_4)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(dff_q_4)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_4)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_4)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_4)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_4)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_4)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(sdpb_inst_113_dout[0]),
  .I1(sdpb_inst_117_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_3)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_3)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_3)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(dff_q_3)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_3)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_3)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(sdpb_inst_105_dout[0]),
  .I1(mux_o_105),
  .S0(dff_q_3)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_106),
  .I1(mux_o_107),
  .S0(dff_q_2)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_110),
  .I1(mux_o_111),
  .S0(dff_q_2)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(dff_q_2)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(dff_q_1)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(dff_q_1)
);
MUX2 mux_inst_120 (
  .O(dout[0]),
  .I0(mux_o_118),
  .I1(mux_o_119),
  .S0(dff_q_0)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(sdpx9b_inst_0_dout[1]),
  .I1(sdpx9b_inst_1_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(sdpx9b_inst_2_dout[1]),
  .I1(sdpx9b_inst_3_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(sdpx9b_inst_4_dout[1]),
  .I1(sdpx9b_inst_5_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(sdpx9b_inst_6_dout[1]),
  .I1(sdpx9b_inst_7_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(sdpx9b_inst_8_dout[1]),
  .I1(sdpx9b_inst_9_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(sdpx9b_inst_10_dout[1]),
  .I1(sdpx9b_inst_11_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(sdpx9b_inst_12_dout[1]),
  .I1(sdpx9b_inst_13_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(sdpx9b_inst_14_dout[1]),
  .I1(sdpx9b_inst_15_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(sdpx9b_inst_16_dout[1]),
  .I1(sdpx9b_inst_17_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(sdpx9b_inst_18_dout[1]),
  .I1(sdpx9b_inst_19_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(sdpx9b_inst_20_dout[1]),
  .I1(sdpx9b_inst_21_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(sdpx9b_inst_22_dout[1]),
  .I1(sdpx9b_inst_23_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(sdpx9b_inst_24_dout[1]),
  .I1(sdpx9b_inst_25_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(sdpx9b_inst_26_dout[1]),
  .I1(sdpx9b_inst_27_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(sdpx9b_inst_28_dout[1]),
  .I1(sdpx9b_inst_29_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(sdpx9b_inst_30_dout[1]),
  .I1(sdpx9b_inst_31_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(sdpx9b_inst_60_dout[1]),
  .I1(sdpx9b_inst_61_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(sdpx9b_inst_62_dout[1]),
  .I1(sdpx9b_inst_63_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(sdpx9b_inst_64_dout[1]),
  .I1(sdpx9b_inst_65_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(sdpx9b_inst_66_dout[1]),
  .I1(sdpx9b_inst_67_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(sdpx9b_inst_68_dout[1]),
  .I1(sdpx9b_inst_69_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(sdpx9b_inst_70_dout[1]),
  .I1(sdpx9b_inst_71_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(sdpx9b_inst_72_dout[1]),
  .I1(sdpx9b_inst_73_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(sdpx9b_inst_74_dout[1]),
  .I1(sdpx9b_inst_75_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(sdpx9b_inst_90_dout[1]),
  .I1(sdpx9b_inst_91_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(sdpx9b_inst_92_dout[1]),
  .I1(sdpx9b_inst_93_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(sdpx9b_inst_94_dout[1]),
  .I1(sdpx9b_inst_95_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(sdpx9b_inst_96_dout[1]),
  .I1(sdpx9b_inst_97_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(dff_q_4)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_4)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_4)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_4)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(dff_q_4)
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(dff_q_4)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(dff_q_4)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(dff_q_4)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_4)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_4)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_4)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_202),
  .I1(mux_o_203),
  .S0(dff_q_4)
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_204),
  .I1(mux_o_205),
  .S0(dff_q_4)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(mux_o_206),
  .I1(mux_o_207),
  .S0(dff_q_4)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(sdpb_inst_113_dout[1]),
  .I1(sdpb_inst_117_dout[1]),
  .S0(dff_q_4)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(mux_o_211),
  .I1(mux_o_212),
  .S0(dff_q_3)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_213),
  .I1(mux_o_214),
  .S0(dff_q_3)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_215),
  .I1(mux_o_216),
  .S0(dff_q_3)
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_3)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_3)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_223),
  .I1(mux_o_224),
  .S0(dff_q_3)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(sdpb_inst_105_dout[1]),
  .I1(mux_o_226),
  .S0(dff_q_3)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(dff_q_2)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(dff_q_2)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_2)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_2)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_1)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_1)
);
MUX2 mux_inst_241 (
  .O(dout[1]),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_0)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(sdpx9b_inst_0_dout[2]),
  .I1(sdpx9b_inst_1_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(sdpx9b_inst_2_dout[2]),
  .I1(sdpx9b_inst_3_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(sdpx9b_inst_4_dout[2]),
  .I1(sdpx9b_inst_5_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(sdpx9b_inst_6_dout[2]),
  .I1(sdpx9b_inst_7_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(sdpx9b_inst_8_dout[2]),
  .I1(sdpx9b_inst_9_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(sdpx9b_inst_10_dout[2]),
  .I1(sdpx9b_inst_11_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(sdpx9b_inst_12_dout[2]),
  .I1(sdpx9b_inst_13_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(sdpx9b_inst_14_dout[2]),
  .I1(sdpx9b_inst_15_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(sdpx9b_inst_16_dout[2]),
  .I1(sdpx9b_inst_17_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(sdpx9b_inst_18_dout[2]),
  .I1(sdpx9b_inst_19_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(sdpx9b_inst_20_dout[2]),
  .I1(sdpx9b_inst_21_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(sdpx9b_inst_22_dout[2]),
  .I1(sdpx9b_inst_23_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(sdpx9b_inst_24_dout[2]),
  .I1(sdpx9b_inst_25_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(sdpx9b_inst_26_dout[2]),
  .I1(sdpx9b_inst_27_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(sdpx9b_inst_28_dout[2]),
  .I1(sdpx9b_inst_29_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(sdpx9b_inst_30_dout[2]),
  .I1(sdpx9b_inst_31_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(sdpx9b_inst_60_dout[2]),
  .I1(sdpx9b_inst_61_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(sdpx9b_inst_62_dout[2]),
  .I1(sdpx9b_inst_63_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(sdpx9b_inst_64_dout[2]),
  .I1(sdpx9b_inst_65_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(sdpx9b_inst_66_dout[2]),
  .I1(sdpx9b_inst_67_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(sdpx9b_inst_68_dout[2]),
  .I1(sdpx9b_inst_69_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(sdpx9b_inst_70_dout[2]),
  .I1(sdpx9b_inst_71_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(sdpx9b_inst_72_dout[2]),
  .I1(sdpx9b_inst_73_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(sdpx9b_inst_74_dout[2]),
  .I1(sdpx9b_inst_75_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(sdpx9b_inst_90_dout[2]),
  .I1(sdpx9b_inst_91_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(sdpx9b_inst_92_dout[2]),
  .I1(sdpx9b_inst_93_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(sdpx9b_inst_94_dout[2]),
  .I1(sdpx9b_inst_95_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(sdpx9b_inst_96_dout[2]),
  .I1(sdpx9b_inst_97_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_4)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_303),
  .I1(mux_o_304),
  .S0(dff_q_4)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_4)
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(mux_o_307),
  .I1(mux_o_308),
  .S0(dff_q_4)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(mux_o_309),
  .I1(mux_o_310),
  .S0(dff_q_4)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(mux_o_311),
  .I1(mux_o_312),
  .S0(dff_q_4)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_313),
  .I1(mux_o_314),
  .S0(dff_q_4)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_4)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_4)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_4)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_321),
  .I1(mux_o_322),
  .S0(dff_q_4)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_323),
  .I1(mux_o_324),
  .S0(dff_q_4)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(mux_o_325),
  .I1(mux_o_326),
  .S0(dff_q_4)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(mux_o_327),
  .I1(mux_o_328),
  .S0(dff_q_4)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(sdpb_inst_113_dout[2]),
  .I1(sdpb_inst_117_dout[2]),
  .S0(dff_q_4)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(dff_q_3)
);
MUX2 mux_inst_349 (
  .O(mux_o_349),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(dff_q_3)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_3)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_3)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_3)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_342),
  .I1(mux_o_343),
  .S0(dff_q_3)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_344),
  .I1(mux_o_345),
  .S0(dff_q_3)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(sdpb_inst_106_dout[2]),
  .I1(mux_o_347),
  .S0(dff_q_3)
);
MUX2 mux_inst_356 (
  .O(mux_o_356),
  .I0(mux_o_348),
  .I1(mux_o_349),
  .S0(dff_q_2)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_2)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_2)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_2)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(mux_o_356),
  .I1(mux_o_357),
  .S0(dff_q_1)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_358),
  .I1(mux_o_359),
  .S0(dff_q_1)
);
MUX2 mux_inst_362 (
  .O(dout[2]),
  .I0(mux_o_360),
  .I1(mux_o_361),
  .S0(dff_q_0)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(sdpx9b_inst_0_dout[3]),
  .I1(sdpx9b_inst_1_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(sdpx9b_inst_2_dout[3]),
  .I1(sdpx9b_inst_3_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(sdpx9b_inst_4_dout[3]),
  .I1(sdpx9b_inst_5_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(sdpx9b_inst_6_dout[3]),
  .I1(sdpx9b_inst_7_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_426 (
  .O(mux_o_426),
  .I0(sdpx9b_inst_8_dout[3]),
  .I1(sdpx9b_inst_9_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(sdpx9b_inst_10_dout[3]),
  .I1(sdpx9b_inst_11_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(sdpx9b_inst_12_dout[3]),
  .I1(sdpx9b_inst_13_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(sdpx9b_inst_14_dout[3]),
  .I1(sdpx9b_inst_15_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(sdpx9b_inst_16_dout[3]),
  .I1(sdpx9b_inst_17_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(sdpx9b_inst_18_dout[3]),
  .I1(sdpx9b_inst_19_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(sdpx9b_inst_20_dout[3]),
  .I1(sdpx9b_inst_21_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_433 (
  .O(mux_o_433),
  .I0(sdpx9b_inst_22_dout[3]),
  .I1(sdpx9b_inst_23_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(sdpx9b_inst_24_dout[3]),
  .I1(sdpx9b_inst_25_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(sdpx9b_inst_26_dout[3]),
  .I1(sdpx9b_inst_27_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(sdpx9b_inst_28_dout[3]),
  .I1(sdpx9b_inst_29_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(sdpx9b_inst_30_dout[3]),
  .I1(sdpx9b_inst_31_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(sdpx9b_inst_60_dout[3]),
  .I1(sdpx9b_inst_61_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(sdpx9b_inst_62_dout[3]),
  .I1(sdpx9b_inst_63_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_440 (
  .O(mux_o_440),
  .I0(sdpx9b_inst_64_dout[3]),
  .I1(sdpx9b_inst_65_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(sdpx9b_inst_66_dout[3]),
  .I1(sdpx9b_inst_67_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(sdpx9b_inst_68_dout[3]),
  .I1(sdpx9b_inst_69_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(sdpx9b_inst_70_dout[3]),
  .I1(sdpx9b_inst_71_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(sdpx9b_inst_72_dout[3]),
  .I1(sdpx9b_inst_73_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(sdpx9b_inst_74_dout[3]),
  .I1(sdpx9b_inst_75_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(sdpx9b_inst_90_dout[3]),
  .I1(sdpx9b_inst_91_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(sdpx9b_inst_92_dout[3]),
  .I1(sdpx9b_inst_93_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(sdpx9b_inst_94_dout[3]),
  .I1(sdpx9b_inst_95_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(sdpx9b_inst_96_dout[3]),
  .I1(sdpx9b_inst_97_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_453 (
  .O(mux_o_453),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(dff_q_4)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(dff_q_4)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_426),
  .I1(mux_o_427),
  .S0(dff_q_4)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_428),
  .I1(mux_o_429),
  .S0(dff_q_4)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_430),
  .I1(mux_o_431),
  .S0(dff_q_4)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_432),
  .I1(mux_o_433),
  .S0(dff_q_4)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(dff_q_4)
);
MUX2 mux_inst_460 (
  .O(mux_o_460),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(dff_q_4)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(dff_q_4)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_440),
  .I1(mux_o_441),
  .S0(dff_q_4)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_442),
  .I1(mux_o_443),
  .S0(dff_q_4)
);
MUX2 mux_inst_464 (
  .O(mux_o_464),
  .I0(mux_o_444),
  .I1(mux_o_445),
  .S0(dff_q_4)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(mux_o_446),
  .I1(mux_o_447),
  .S0(dff_q_4)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(mux_o_448),
  .I1(mux_o_449),
  .S0(dff_q_4)
);
MUX2 mux_inst_468 (
  .O(mux_o_468),
  .I0(sdpb_inst_113_dout[3]),
  .I1(sdpb_inst_117_dout[3]),
  .S0(dff_q_4)
);
MUX2 mux_inst_469 (
  .O(mux_o_469),
  .I0(mux_o_453),
  .I1(mux_o_454),
  .S0(dff_q_3)
);
MUX2 mux_inst_470 (
  .O(mux_o_470),
  .I0(mux_o_455),
  .I1(mux_o_456),
  .S0(dff_q_3)
);
MUX2 mux_inst_471 (
  .O(mux_o_471),
  .I0(mux_o_457),
  .I1(mux_o_458),
  .S0(dff_q_3)
);
MUX2 mux_inst_472 (
  .O(mux_o_472),
  .I0(mux_o_459),
  .I1(mux_o_460),
  .S0(dff_q_3)
);
MUX2 mux_inst_473 (
  .O(mux_o_473),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(dff_q_3)
);
MUX2 mux_inst_474 (
  .O(mux_o_474),
  .I0(mux_o_463),
  .I1(mux_o_464),
  .S0(dff_q_3)
);
MUX2 mux_inst_475 (
  .O(mux_o_475),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_3)
);
MUX2 mux_inst_476 (
  .O(mux_o_476),
  .I0(sdpb_inst_106_dout[3]),
  .I1(mux_o_468),
  .S0(dff_q_3)
);
MUX2 mux_inst_477 (
  .O(mux_o_477),
  .I0(mux_o_469),
  .I1(mux_o_470),
  .S0(dff_q_2)
);
MUX2 mux_inst_478 (
  .O(mux_o_478),
  .I0(mux_o_471),
  .I1(mux_o_472),
  .S0(dff_q_2)
);
MUX2 mux_inst_479 (
  .O(mux_o_479),
  .I0(mux_o_473),
  .I1(mux_o_474),
  .S0(dff_q_2)
);
MUX2 mux_inst_480 (
  .O(mux_o_480),
  .I0(mux_o_475),
  .I1(mux_o_476),
  .S0(dff_q_2)
);
MUX2 mux_inst_481 (
  .O(mux_o_481),
  .I0(mux_o_477),
  .I1(mux_o_478),
  .S0(dff_q_1)
);
MUX2 mux_inst_482 (
  .O(mux_o_482),
  .I0(mux_o_479),
  .I1(mux_o_480),
  .S0(dff_q_1)
);
MUX2 mux_inst_483 (
  .O(dout[3]),
  .I0(mux_o_481),
  .I1(mux_o_482),
  .S0(dff_q_0)
);
MUX2 mux_inst_543 (
  .O(mux_o_543),
  .I0(sdpx9b_inst_0_dout[4]),
  .I1(sdpx9b_inst_1_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_544 (
  .O(mux_o_544),
  .I0(sdpx9b_inst_2_dout[4]),
  .I1(sdpx9b_inst_3_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_545 (
  .O(mux_o_545),
  .I0(sdpx9b_inst_4_dout[4]),
  .I1(sdpx9b_inst_5_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_546 (
  .O(mux_o_546),
  .I0(sdpx9b_inst_6_dout[4]),
  .I1(sdpx9b_inst_7_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_547 (
  .O(mux_o_547),
  .I0(sdpx9b_inst_8_dout[4]),
  .I1(sdpx9b_inst_9_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_548 (
  .O(mux_o_548),
  .I0(sdpx9b_inst_10_dout[4]),
  .I1(sdpx9b_inst_11_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_549 (
  .O(mux_o_549),
  .I0(sdpx9b_inst_12_dout[4]),
  .I1(sdpx9b_inst_13_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_550 (
  .O(mux_o_550),
  .I0(sdpx9b_inst_14_dout[4]),
  .I1(sdpx9b_inst_15_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_551 (
  .O(mux_o_551),
  .I0(sdpx9b_inst_16_dout[4]),
  .I1(sdpx9b_inst_17_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_552 (
  .O(mux_o_552),
  .I0(sdpx9b_inst_18_dout[4]),
  .I1(sdpx9b_inst_19_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_553 (
  .O(mux_o_553),
  .I0(sdpx9b_inst_20_dout[4]),
  .I1(sdpx9b_inst_21_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_554 (
  .O(mux_o_554),
  .I0(sdpx9b_inst_22_dout[4]),
  .I1(sdpx9b_inst_23_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_555 (
  .O(mux_o_555),
  .I0(sdpx9b_inst_24_dout[4]),
  .I1(sdpx9b_inst_25_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_556 (
  .O(mux_o_556),
  .I0(sdpx9b_inst_26_dout[4]),
  .I1(sdpx9b_inst_27_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_557 (
  .O(mux_o_557),
  .I0(sdpx9b_inst_28_dout[4]),
  .I1(sdpx9b_inst_29_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_558 (
  .O(mux_o_558),
  .I0(sdpx9b_inst_30_dout[4]),
  .I1(sdpx9b_inst_31_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_559 (
  .O(mux_o_559),
  .I0(sdpx9b_inst_60_dout[4]),
  .I1(sdpx9b_inst_61_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(sdpx9b_inst_62_dout[4]),
  .I1(sdpx9b_inst_63_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(sdpx9b_inst_64_dout[4]),
  .I1(sdpx9b_inst_65_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_562 (
  .O(mux_o_562),
  .I0(sdpx9b_inst_66_dout[4]),
  .I1(sdpx9b_inst_67_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_563 (
  .O(mux_o_563),
  .I0(sdpx9b_inst_68_dout[4]),
  .I1(sdpx9b_inst_69_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_564 (
  .O(mux_o_564),
  .I0(sdpx9b_inst_70_dout[4]),
  .I1(sdpx9b_inst_71_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_565 (
  .O(mux_o_565),
  .I0(sdpx9b_inst_72_dout[4]),
  .I1(sdpx9b_inst_73_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_566 (
  .O(mux_o_566),
  .I0(sdpx9b_inst_74_dout[4]),
  .I1(sdpx9b_inst_75_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_567 (
  .O(mux_o_567),
  .I0(sdpx9b_inst_90_dout[4]),
  .I1(sdpx9b_inst_91_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_568 (
  .O(mux_o_568),
  .I0(sdpx9b_inst_92_dout[4]),
  .I1(sdpx9b_inst_93_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_569 (
  .O(mux_o_569),
  .I0(sdpx9b_inst_94_dout[4]),
  .I1(sdpx9b_inst_95_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_570 (
  .O(mux_o_570),
  .I0(sdpx9b_inst_96_dout[4]),
  .I1(sdpx9b_inst_97_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_574 (
  .O(mux_o_574),
  .I0(mux_o_543),
  .I1(mux_o_544),
  .S0(dff_q_4)
);
MUX2 mux_inst_575 (
  .O(mux_o_575),
  .I0(mux_o_545),
  .I1(mux_o_546),
  .S0(dff_q_4)
);
MUX2 mux_inst_576 (
  .O(mux_o_576),
  .I0(mux_o_547),
  .I1(mux_o_548),
  .S0(dff_q_4)
);
MUX2 mux_inst_577 (
  .O(mux_o_577),
  .I0(mux_o_549),
  .I1(mux_o_550),
  .S0(dff_q_4)
);
MUX2 mux_inst_578 (
  .O(mux_o_578),
  .I0(mux_o_551),
  .I1(mux_o_552),
  .S0(dff_q_4)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(mux_o_553),
  .I1(mux_o_554),
  .S0(dff_q_4)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(mux_o_555),
  .I1(mux_o_556),
  .S0(dff_q_4)
);
MUX2 mux_inst_581 (
  .O(mux_o_581),
  .I0(mux_o_557),
  .I1(mux_o_558),
  .S0(dff_q_4)
);
MUX2 mux_inst_582 (
  .O(mux_o_582),
  .I0(mux_o_559),
  .I1(mux_o_560),
  .S0(dff_q_4)
);
MUX2 mux_inst_583 (
  .O(mux_o_583),
  .I0(mux_o_561),
  .I1(mux_o_562),
  .S0(dff_q_4)
);
MUX2 mux_inst_584 (
  .O(mux_o_584),
  .I0(mux_o_563),
  .I1(mux_o_564),
  .S0(dff_q_4)
);
MUX2 mux_inst_585 (
  .O(mux_o_585),
  .I0(mux_o_565),
  .I1(mux_o_566),
  .S0(dff_q_4)
);
MUX2 mux_inst_586 (
  .O(mux_o_586),
  .I0(mux_o_567),
  .I1(mux_o_568),
  .S0(dff_q_4)
);
MUX2 mux_inst_587 (
  .O(mux_o_587),
  .I0(mux_o_569),
  .I1(mux_o_570),
  .S0(dff_q_4)
);
MUX2 mux_inst_589 (
  .O(mux_o_589),
  .I0(sdpb_inst_114_dout[4]),
  .I1(sdpb_inst_117_dout[4]),
  .S0(dff_q_4)
);
MUX2 mux_inst_590 (
  .O(mux_o_590),
  .I0(mux_o_574),
  .I1(mux_o_575),
  .S0(dff_q_3)
);
MUX2 mux_inst_591 (
  .O(mux_o_591),
  .I0(mux_o_576),
  .I1(mux_o_577),
  .S0(dff_q_3)
);
MUX2 mux_inst_592 (
  .O(mux_o_592),
  .I0(mux_o_578),
  .I1(mux_o_579),
  .S0(dff_q_3)
);
MUX2 mux_inst_593 (
  .O(mux_o_593),
  .I0(mux_o_580),
  .I1(mux_o_581),
  .S0(dff_q_3)
);
MUX2 mux_inst_594 (
  .O(mux_o_594),
  .I0(mux_o_582),
  .I1(mux_o_583),
  .S0(dff_q_3)
);
MUX2 mux_inst_595 (
  .O(mux_o_595),
  .I0(mux_o_584),
  .I1(mux_o_585),
  .S0(dff_q_3)
);
MUX2 mux_inst_596 (
  .O(mux_o_596),
  .I0(mux_o_586),
  .I1(mux_o_587),
  .S0(dff_q_3)
);
MUX2 mux_inst_597 (
  .O(mux_o_597),
  .I0(sdpb_inst_107_dout[4]),
  .I1(mux_o_589),
  .S0(dff_q_3)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(mux_o_590),
  .I1(mux_o_591),
  .S0(dff_q_2)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(mux_o_592),
  .I1(mux_o_593),
  .S0(dff_q_2)
);
MUX2 mux_inst_600 (
  .O(mux_o_600),
  .I0(mux_o_594),
  .I1(mux_o_595),
  .S0(dff_q_2)
);
MUX2 mux_inst_601 (
  .O(mux_o_601),
  .I0(mux_o_596),
  .I1(mux_o_597),
  .S0(dff_q_2)
);
MUX2 mux_inst_602 (
  .O(mux_o_602),
  .I0(mux_o_598),
  .I1(mux_o_599),
  .S0(dff_q_1)
);
MUX2 mux_inst_603 (
  .O(mux_o_603),
  .I0(mux_o_600),
  .I1(mux_o_601),
  .S0(dff_q_1)
);
MUX2 mux_inst_604 (
  .O(dout[4]),
  .I0(mux_o_602),
  .I1(mux_o_603),
  .S0(dff_q_0)
);
MUX2 mux_inst_664 (
  .O(mux_o_664),
  .I0(sdpx9b_inst_0_dout[5]),
  .I1(sdpx9b_inst_1_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_665 (
  .O(mux_o_665),
  .I0(sdpx9b_inst_2_dout[5]),
  .I1(sdpx9b_inst_3_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_666 (
  .O(mux_o_666),
  .I0(sdpx9b_inst_4_dout[5]),
  .I1(sdpx9b_inst_5_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_667 (
  .O(mux_o_667),
  .I0(sdpx9b_inst_6_dout[5]),
  .I1(sdpx9b_inst_7_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_668 (
  .O(mux_o_668),
  .I0(sdpx9b_inst_8_dout[5]),
  .I1(sdpx9b_inst_9_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_669 (
  .O(mux_o_669),
  .I0(sdpx9b_inst_10_dout[5]),
  .I1(sdpx9b_inst_11_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_670 (
  .O(mux_o_670),
  .I0(sdpx9b_inst_12_dout[5]),
  .I1(sdpx9b_inst_13_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_671 (
  .O(mux_o_671),
  .I0(sdpx9b_inst_14_dout[5]),
  .I1(sdpx9b_inst_15_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_672 (
  .O(mux_o_672),
  .I0(sdpx9b_inst_16_dout[5]),
  .I1(sdpx9b_inst_17_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_673 (
  .O(mux_o_673),
  .I0(sdpx9b_inst_18_dout[5]),
  .I1(sdpx9b_inst_19_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_674 (
  .O(mux_o_674),
  .I0(sdpx9b_inst_20_dout[5]),
  .I1(sdpx9b_inst_21_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_675 (
  .O(mux_o_675),
  .I0(sdpx9b_inst_22_dout[5]),
  .I1(sdpx9b_inst_23_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_676 (
  .O(mux_o_676),
  .I0(sdpx9b_inst_24_dout[5]),
  .I1(sdpx9b_inst_25_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_677 (
  .O(mux_o_677),
  .I0(sdpx9b_inst_26_dout[5]),
  .I1(sdpx9b_inst_27_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_678 (
  .O(mux_o_678),
  .I0(sdpx9b_inst_28_dout[5]),
  .I1(sdpx9b_inst_29_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_679 (
  .O(mux_o_679),
  .I0(sdpx9b_inst_30_dout[5]),
  .I1(sdpx9b_inst_31_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_680 (
  .O(mux_o_680),
  .I0(sdpx9b_inst_60_dout[5]),
  .I1(sdpx9b_inst_61_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_681 (
  .O(mux_o_681),
  .I0(sdpx9b_inst_62_dout[5]),
  .I1(sdpx9b_inst_63_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_682 (
  .O(mux_o_682),
  .I0(sdpx9b_inst_64_dout[5]),
  .I1(sdpx9b_inst_65_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_683 (
  .O(mux_o_683),
  .I0(sdpx9b_inst_66_dout[5]),
  .I1(sdpx9b_inst_67_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_684 (
  .O(mux_o_684),
  .I0(sdpx9b_inst_68_dout[5]),
  .I1(sdpx9b_inst_69_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_685 (
  .O(mux_o_685),
  .I0(sdpx9b_inst_70_dout[5]),
  .I1(sdpx9b_inst_71_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_686 (
  .O(mux_o_686),
  .I0(sdpx9b_inst_72_dout[5]),
  .I1(sdpx9b_inst_73_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_687 (
  .O(mux_o_687),
  .I0(sdpx9b_inst_74_dout[5]),
  .I1(sdpx9b_inst_75_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_688 (
  .O(mux_o_688),
  .I0(sdpx9b_inst_90_dout[5]),
  .I1(sdpx9b_inst_91_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_689 (
  .O(mux_o_689),
  .I0(sdpx9b_inst_92_dout[5]),
  .I1(sdpx9b_inst_93_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_690 (
  .O(mux_o_690),
  .I0(sdpx9b_inst_94_dout[5]),
  .I1(sdpx9b_inst_95_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_691 (
  .O(mux_o_691),
  .I0(sdpx9b_inst_96_dout[5]),
  .I1(sdpx9b_inst_97_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_695 (
  .O(mux_o_695),
  .I0(mux_o_664),
  .I1(mux_o_665),
  .S0(dff_q_4)
);
MUX2 mux_inst_696 (
  .O(mux_o_696),
  .I0(mux_o_666),
  .I1(mux_o_667),
  .S0(dff_q_4)
);
MUX2 mux_inst_697 (
  .O(mux_o_697),
  .I0(mux_o_668),
  .I1(mux_o_669),
  .S0(dff_q_4)
);
MUX2 mux_inst_698 (
  .O(mux_o_698),
  .I0(mux_o_670),
  .I1(mux_o_671),
  .S0(dff_q_4)
);
MUX2 mux_inst_699 (
  .O(mux_o_699),
  .I0(mux_o_672),
  .I1(mux_o_673),
  .S0(dff_q_4)
);
MUX2 mux_inst_700 (
  .O(mux_o_700),
  .I0(mux_o_674),
  .I1(mux_o_675),
  .S0(dff_q_4)
);
MUX2 mux_inst_701 (
  .O(mux_o_701),
  .I0(mux_o_676),
  .I1(mux_o_677),
  .S0(dff_q_4)
);
MUX2 mux_inst_702 (
  .O(mux_o_702),
  .I0(mux_o_678),
  .I1(mux_o_679),
  .S0(dff_q_4)
);
MUX2 mux_inst_703 (
  .O(mux_o_703),
  .I0(mux_o_680),
  .I1(mux_o_681),
  .S0(dff_q_4)
);
MUX2 mux_inst_704 (
  .O(mux_o_704),
  .I0(mux_o_682),
  .I1(mux_o_683),
  .S0(dff_q_4)
);
MUX2 mux_inst_705 (
  .O(mux_o_705),
  .I0(mux_o_684),
  .I1(mux_o_685),
  .S0(dff_q_4)
);
MUX2 mux_inst_706 (
  .O(mux_o_706),
  .I0(mux_o_686),
  .I1(mux_o_687),
  .S0(dff_q_4)
);
MUX2 mux_inst_707 (
  .O(mux_o_707),
  .I0(mux_o_688),
  .I1(mux_o_689),
  .S0(dff_q_4)
);
MUX2 mux_inst_708 (
  .O(mux_o_708),
  .I0(mux_o_690),
  .I1(mux_o_691),
  .S0(dff_q_4)
);
MUX2 mux_inst_710 (
  .O(mux_o_710),
  .I0(sdpb_inst_114_dout[5]),
  .I1(sdpb_inst_117_dout[5]),
  .S0(dff_q_4)
);
MUX2 mux_inst_711 (
  .O(mux_o_711),
  .I0(mux_o_695),
  .I1(mux_o_696),
  .S0(dff_q_3)
);
MUX2 mux_inst_712 (
  .O(mux_o_712),
  .I0(mux_o_697),
  .I1(mux_o_698),
  .S0(dff_q_3)
);
MUX2 mux_inst_713 (
  .O(mux_o_713),
  .I0(mux_o_699),
  .I1(mux_o_700),
  .S0(dff_q_3)
);
MUX2 mux_inst_714 (
  .O(mux_o_714),
  .I0(mux_o_701),
  .I1(mux_o_702),
  .S0(dff_q_3)
);
MUX2 mux_inst_715 (
  .O(mux_o_715),
  .I0(mux_o_703),
  .I1(mux_o_704),
  .S0(dff_q_3)
);
MUX2 mux_inst_716 (
  .O(mux_o_716),
  .I0(mux_o_705),
  .I1(mux_o_706),
  .S0(dff_q_3)
);
MUX2 mux_inst_717 (
  .O(mux_o_717),
  .I0(mux_o_707),
  .I1(mux_o_708),
  .S0(dff_q_3)
);
MUX2 mux_inst_718 (
  .O(mux_o_718),
  .I0(sdpb_inst_107_dout[5]),
  .I1(mux_o_710),
  .S0(dff_q_3)
);
MUX2 mux_inst_719 (
  .O(mux_o_719),
  .I0(mux_o_711),
  .I1(mux_o_712),
  .S0(dff_q_2)
);
MUX2 mux_inst_720 (
  .O(mux_o_720),
  .I0(mux_o_713),
  .I1(mux_o_714),
  .S0(dff_q_2)
);
MUX2 mux_inst_721 (
  .O(mux_o_721),
  .I0(mux_o_715),
  .I1(mux_o_716),
  .S0(dff_q_2)
);
MUX2 mux_inst_722 (
  .O(mux_o_722),
  .I0(mux_o_717),
  .I1(mux_o_718),
  .S0(dff_q_2)
);
MUX2 mux_inst_723 (
  .O(mux_o_723),
  .I0(mux_o_719),
  .I1(mux_o_720),
  .S0(dff_q_1)
);
MUX2 mux_inst_724 (
  .O(mux_o_724),
  .I0(mux_o_721),
  .I1(mux_o_722),
  .S0(dff_q_1)
);
MUX2 mux_inst_725 (
  .O(dout[5]),
  .I0(mux_o_723),
  .I1(mux_o_724),
  .S0(dff_q_0)
);
MUX2 mux_inst_785 (
  .O(mux_o_785),
  .I0(sdpx9b_inst_0_dout[6]),
  .I1(sdpx9b_inst_1_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_786 (
  .O(mux_o_786),
  .I0(sdpx9b_inst_2_dout[6]),
  .I1(sdpx9b_inst_3_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_787 (
  .O(mux_o_787),
  .I0(sdpx9b_inst_4_dout[6]),
  .I1(sdpx9b_inst_5_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_788 (
  .O(mux_o_788),
  .I0(sdpx9b_inst_6_dout[6]),
  .I1(sdpx9b_inst_7_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_789 (
  .O(mux_o_789),
  .I0(sdpx9b_inst_8_dout[6]),
  .I1(sdpx9b_inst_9_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_790 (
  .O(mux_o_790),
  .I0(sdpx9b_inst_10_dout[6]),
  .I1(sdpx9b_inst_11_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_791 (
  .O(mux_o_791),
  .I0(sdpx9b_inst_12_dout[6]),
  .I1(sdpx9b_inst_13_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_792 (
  .O(mux_o_792),
  .I0(sdpx9b_inst_14_dout[6]),
  .I1(sdpx9b_inst_15_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_793 (
  .O(mux_o_793),
  .I0(sdpx9b_inst_16_dout[6]),
  .I1(sdpx9b_inst_17_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_794 (
  .O(mux_o_794),
  .I0(sdpx9b_inst_18_dout[6]),
  .I1(sdpx9b_inst_19_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_795 (
  .O(mux_o_795),
  .I0(sdpx9b_inst_20_dout[6]),
  .I1(sdpx9b_inst_21_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_796 (
  .O(mux_o_796),
  .I0(sdpx9b_inst_22_dout[6]),
  .I1(sdpx9b_inst_23_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_797 (
  .O(mux_o_797),
  .I0(sdpx9b_inst_24_dout[6]),
  .I1(sdpx9b_inst_25_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_798 (
  .O(mux_o_798),
  .I0(sdpx9b_inst_26_dout[6]),
  .I1(sdpx9b_inst_27_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_799 (
  .O(mux_o_799),
  .I0(sdpx9b_inst_28_dout[6]),
  .I1(sdpx9b_inst_29_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_800 (
  .O(mux_o_800),
  .I0(sdpx9b_inst_30_dout[6]),
  .I1(sdpx9b_inst_31_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_801 (
  .O(mux_o_801),
  .I0(sdpx9b_inst_60_dout[6]),
  .I1(sdpx9b_inst_61_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_802 (
  .O(mux_o_802),
  .I0(sdpx9b_inst_62_dout[6]),
  .I1(sdpx9b_inst_63_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_803 (
  .O(mux_o_803),
  .I0(sdpx9b_inst_64_dout[6]),
  .I1(sdpx9b_inst_65_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_804 (
  .O(mux_o_804),
  .I0(sdpx9b_inst_66_dout[6]),
  .I1(sdpx9b_inst_67_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_805 (
  .O(mux_o_805),
  .I0(sdpx9b_inst_68_dout[6]),
  .I1(sdpx9b_inst_69_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_806 (
  .O(mux_o_806),
  .I0(sdpx9b_inst_70_dout[6]),
  .I1(sdpx9b_inst_71_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_807 (
  .O(mux_o_807),
  .I0(sdpx9b_inst_72_dout[6]),
  .I1(sdpx9b_inst_73_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_808 (
  .O(mux_o_808),
  .I0(sdpx9b_inst_74_dout[6]),
  .I1(sdpx9b_inst_75_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_809 (
  .O(mux_o_809),
  .I0(sdpx9b_inst_90_dout[6]),
  .I1(sdpx9b_inst_91_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_810 (
  .O(mux_o_810),
  .I0(sdpx9b_inst_92_dout[6]),
  .I1(sdpx9b_inst_93_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_811 (
  .O(mux_o_811),
  .I0(sdpx9b_inst_94_dout[6]),
  .I1(sdpx9b_inst_95_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_812 (
  .O(mux_o_812),
  .I0(sdpx9b_inst_96_dout[6]),
  .I1(sdpx9b_inst_97_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_816 (
  .O(mux_o_816),
  .I0(mux_o_785),
  .I1(mux_o_786),
  .S0(dff_q_4)
);
MUX2 mux_inst_817 (
  .O(mux_o_817),
  .I0(mux_o_787),
  .I1(mux_o_788),
  .S0(dff_q_4)
);
MUX2 mux_inst_818 (
  .O(mux_o_818),
  .I0(mux_o_789),
  .I1(mux_o_790),
  .S0(dff_q_4)
);
MUX2 mux_inst_819 (
  .O(mux_o_819),
  .I0(mux_o_791),
  .I1(mux_o_792),
  .S0(dff_q_4)
);
MUX2 mux_inst_820 (
  .O(mux_o_820),
  .I0(mux_o_793),
  .I1(mux_o_794),
  .S0(dff_q_4)
);
MUX2 mux_inst_821 (
  .O(mux_o_821),
  .I0(mux_o_795),
  .I1(mux_o_796),
  .S0(dff_q_4)
);
MUX2 mux_inst_822 (
  .O(mux_o_822),
  .I0(mux_o_797),
  .I1(mux_o_798),
  .S0(dff_q_4)
);
MUX2 mux_inst_823 (
  .O(mux_o_823),
  .I0(mux_o_799),
  .I1(mux_o_800),
  .S0(dff_q_4)
);
MUX2 mux_inst_824 (
  .O(mux_o_824),
  .I0(mux_o_801),
  .I1(mux_o_802),
  .S0(dff_q_4)
);
MUX2 mux_inst_825 (
  .O(mux_o_825),
  .I0(mux_o_803),
  .I1(mux_o_804),
  .S0(dff_q_4)
);
MUX2 mux_inst_826 (
  .O(mux_o_826),
  .I0(mux_o_805),
  .I1(mux_o_806),
  .S0(dff_q_4)
);
MUX2 mux_inst_827 (
  .O(mux_o_827),
  .I0(mux_o_807),
  .I1(mux_o_808),
  .S0(dff_q_4)
);
MUX2 mux_inst_828 (
  .O(mux_o_828),
  .I0(mux_o_809),
  .I1(mux_o_810),
  .S0(dff_q_4)
);
MUX2 mux_inst_829 (
  .O(mux_o_829),
  .I0(mux_o_811),
  .I1(mux_o_812),
  .S0(dff_q_4)
);
MUX2 mux_inst_831 (
  .O(mux_o_831),
  .I0(sdpb_inst_114_dout[6]),
  .I1(sdpb_inst_117_dout[6]),
  .S0(dff_q_4)
);
MUX2 mux_inst_832 (
  .O(mux_o_832),
  .I0(mux_o_816),
  .I1(mux_o_817),
  .S0(dff_q_3)
);
MUX2 mux_inst_833 (
  .O(mux_o_833),
  .I0(mux_o_818),
  .I1(mux_o_819),
  .S0(dff_q_3)
);
MUX2 mux_inst_834 (
  .O(mux_o_834),
  .I0(mux_o_820),
  .I1(mux_o_821),
  .S0(dff_q_3)
);
MUX2 mux_inst_835 (
  .O(mux_o_835),
  .I0(mux_o_822),
  .I1(mux_o_823),
  .S0(dff_q_3)
);
MUX2 mux_inst_836 (
  .O(mux_o_836),
  .I0(mux_o_824),
  .I1(mux_o_825),
  .S0(dff_q_3)
);
MUX2 mux_inst_837 (
  .O(mux_o_837),
  .I0(mux_o_826),
  .I1(mux_o_827),
  .S0(dff_q_3)
);
MUX2 mux_inst_838 (
  .O(mux_o_838),
  .I0(mux_o_828),
  .I1(mux_o_829),
  .S0(dff_q_3)
);
MUX2 mux_inst_839 (
  .O(mux_o_839),
  .I0(sdpb_inst_108_dout[6]),
  .I1(mux_o_831),
  .S0(dff_q_3)
);
MUX2 mux_inst_840 (
  .O(mux_o_840),
  .I0(mux_o_832),
  .I1(mux_o_833),
  .S0(dff_q_2)
);
MUX2 mux_inst_841 (
  .O(mux_o_841),
  .I0(mux_o_834),
  .I1(mux_o_835),
  .S0(dff_q_2)
);
MUX2 mux_inst_842 (
  .O(mux_o_842),
  .I0(mux_o_836),
  .I1(mux_o_837),
  .S0(dff_q_2)
);
MUX2 mux_inst_843 (
  .O(mux_o_843),
  .I0(mux_o_838),
  .I1(mux_o_839),
  .S0(dff_q_2)
);
MUX2 mux_inst_844 (
  .O(mux_o_844),
  .I0(mux_o_840),
  .I1(mux_o_841),
  .S0(dff_q_1)
);
MUX2 mux_inst_845 (
  .O(mux_o_845),
  .I0(mux_o_842),
  .I1(mux_o_843),
  .S0(dff_q_1)
);
MUX2 mux_inst_846 (
  .O(dout[6]),
  .I0(mux_o_844),
  .I1(mux_o_845),
  .S0(dff_q_0)
);
MUX2 mux_inst_906 (
  .O(mux_o_906),
  .I0(sdpx9b_inst_0_dout[7]),
  .I1(sdpx9b_inst_1_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_907 (
  .O(mux_o_907),
  .I0(sdpx9b_inst_2_dout[7]),
  .I1(sdpx9b_inst_3_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_908 (
  .O(mux_o_908),
  .I0(sdpx9b_inst_4_dout[7]),
  .I1(sdpx9b_inst_5_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_909 (
  .O(mux_o_909),
  .I0(sdpx9b_inst_6_dout[7]),
  .I1(sdpx9b_inst_7_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_910 (
  .O(mux_o_910),
  .I0(sdpx9b_inst_8_dout[7]),
  .I1(sdpx9b_inst_9_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_911 (
  .O(mux_o_911),
  .I0(sdpx9b_inst_10_dout[7]),
  .I1(sdpx9b_inst_11_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_912 (
  .O(mux_o_912),
  .I0(sdpx9b_inst_12_dout[7]),
  .I1(sdpx9b_inst_13_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_913 (
  .O(mux_o_913),
  .I0(sdpx9b_inst_14_dout[7]),
  .I1(sdpx9b_inst_15_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_914 (
  .O(mux_o_914),
  .I0(sdpx9b_inst_16_dout[7]),
  .I1(sdpx9b_inst_17_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_915 (
  .O(mux_o_915),
  .I0(sdpx9b_inst_18_dout[7]),
  .I1(sdpx9b_inst_19_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_916 (
  .O(mux_o_916),
  .I0(sdpx9b_inst_20_dout[7]),
  .I1(sdpx9b_inst_21_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_917 (
  .O(mux_o_917),
  .I0(sdpx9b_inst_22_dout[7]),
  .I1(sdpx9b_inst_23_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_918 (
  .O(mux_o_918),
  .I0(sdpx9b_inst_24_dout[7]),
  .I1(sdpx9b_inst_25_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_919 (
  .O(mux_o_919),
  .I0(sdpx9b_inst_26_dout[7]),
  .I1(sdpx9b_inst_27_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_920 (
  .O(mux_o_920),
  .I0(sdpx9b_inst_28_dout[7]),
  .I1(sdpx9b_inst_29_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_921 (
  .O(mux_o_921),
  .I0(sdpx9b_inst_30_dout[7]),
  .I1(sdpx9b_inst_31_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_922 (
  .O(mux_o_922),
  .I0(sdpx9b_inst_60_dout[7]),
  .I1(sdpx9b_inst_61_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_923 (
  .O(mux_o_923),
  .I0(sdpx9b_inst_62_dout[7]),
  .I1(sdpx9b_inst_63_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_924 (
  .O(mux_o_924),
  .I0(sdpx9b_inst_64_dout[7]),
  .I1(sdpx9b_inst_65_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_925 (
  .O(mux_o_925),
  .I0(sdpx9b_inst_66_dout[7]),
  .I1(sdpx9b_inst_67_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_926 (
  .O(mux_o_926),
  .I0(sdpx9b_inst_68_dout[7]),
  .I1(sdpx9b_inst_69_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_927 (
  .O(mux_o_927),
  .I0(sdpx9b_inst_70_dout[7]),
  .I1(sdpx9b_inst_71_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_928 (
  .O(mux_o_928),
  .I0(sdpx9b_inst_72_dout[7]),
  .I1(sdpx9b_inst_73_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_929 (
  .O(mux_o_929),
  .I0(sdpx9b_inst_74_dout[7]),
  .I1(sdpx9b_inst_75_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_930 (
  .O(mux_o_930),
  .I0(sdpx9b_inst_90_dout[7]),
  .I1(sdpx9b_inst_91_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_931 (
  .O(mux_o_931),
  .I0(sdpx9b_inst_92_dout[7]),
  .I1(sdpx9b_inst_93_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_932 (
  .O(mux_o_932),
  .I0(sdpx9b_inst_94_dout[7]),
  .I1(sdpx9b_inst_95_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_933 (
  .O(mux_o_933),
  .I0(sdpx9b_inst_96_dout[7]),
  .I1(sdpx9b_inst_97_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_937 (
  .O(mux_o_937),
  .I0(mux_o_906),
  .I1(mux_o_907),
  .S0(dff_q_4)
);
MUX2 mux_inst_938 (
  .O(mux_o_938),
  .I0(mux_o_908),
  .I1(mux_o_909),
  .S0(dff_q_4)
);
MUX2 mux_inst_939 (
  .O(mux_o_939),
  .I0(mux_o_910),
  .I1(mux_o_911),
  .S0(dff_q_4)
);
MUX2 mux_inst_940 (
  .O(mux_o_940),
  .I0(mux_o_912),
  .I1(mux_o_913),
  .S0(dff_q_4)
);
MUX2 mux_inst_941 (
  .O(mux_o_941),
  .I0(mux_o_914),
  .I1(mux_o_915),
  .S0(dff_q_4)
);
MUX2 mux_inst_942 (
  .O(mux_o_942),
  .I0(mux_o_916),
  .I1(mux_o_917),
  .S0(dff_q_4)
);
MUX2 mux_inst_943 (
  .O(mux_o_943),
  .I0(mux_o_918),
  .I1(mux_o_919),
  .S0(dff_q_4)
);
MUX2 mux_inst_944 (
  .O(mux_o_944),
  .I0(mux_o_920),
  .I1(mux_o_921),
  .S0(dff_q_4)
);
MUX2 mux_inst_945 (
  .O(mux_o_945),
  .I0(mux_o_922),
  .I1(mux_o_923),
  .S0(dff_q_4)
);
MUX2 mux_inst_946 (
  .O(mux_o_946),
  .I0(mux_o_924),
  .I1(mux_o_925),
  .S0(dff_q_4)
);
MUX2 mux_inst_947 (
  .O(mux_o_947),
  .I0(mux_o_926),
  .I1(mux_o_927),
  .S0(dff_q_4)
);
MUX2 mux_inst_948 (
  .O(mux_o_948),
  .I0(mux_o_928),
  .I1(mux_o_929),
  .S0(dff_q_4)
);
MUX2 mux_inst_949 (
  .O(mux_o_949),
  .I0(mux_o_930),
  .I1(mux_o_931),
  .S0(dff_q_4)
);
MUX2 mux_inst_950 (
  .O(mux_o_950),
  .I0(mux_o_932),
  .I1(mux_o_933),
  .S0(dff_q_4)
);
MUX2 mux_inst_952 (
  .O(mux_o_952),
  .I0(sdpb_inst_114_dout[7]),
  .I1(sdpb_inst_117_dout[7]),
  .S0(dff_q_4)
);
MUX2 mux_inst_953 (
  .O(mux_o_953),
  .I0(mux_o_937),
  .I1(mux_o_938),
  .S0(dff_q_3)
);
MUX2 mux_inst_954 (
  .O(mux_o_954),
  .I0(mux_o_939),
  .I1(mux_o_940),
  .S0(dff_q_3)
);
MUX2 mux_inst_955 (
  .O(mux_o_955),
  .I0(mux_o_941),
  .I1(mux_o_942),
  .S0(dff_q_3)
);
MUX2 mux_inst_956 (
  .O(mux_o_956),
  .I0(mux_o_943),
  .I1(mux_o_944),
  .S0(dff_q_3)
);
MUX2 mux_inst_957 (
  .O(mux_o_957),
  .I0(mux_o_945),
  .I1(mux_o_946),
  .S0(dff_q_3)
);
MUX2 mux_inst_958 (
  .O(mux_o_958),
  .I0(mux_o_947),
  .I1(mux_o_948),
  .S0(dff_q_3)
);
MUX2 mux_inst_959 (
  .O(mux_o_959),
  .I0(mux_o_949),
  .I1(mux_o_950),
  .S0(dff_q_3)
);
MUX2 mux_inst_960 (
  .O(mux_o_960),
  .I0(sdpb_inst_108_dout[7]),
  .I1(mux_o_952),
  .S0(dff_q_3)
);
MUX2 mux_inst_961 (
  .O(mux_o_961),
  .I0(mux_o_953),
  .I1(mux_o_954),
  .S0(dff_q_2)
);
MUX2 mux_inst_962 (
  .O(mux_o_962),
  .I0(mux_o_955),
  .I1(mux_o_956),
  .S0(dff_q_2)
);
MUX2 mux_inst_963 (
  .O(mux_o_963),
  .I0(mux_o_957),
  .I1(mux_o_958),
  .S0(dff_q_2)
);
MUX2 mux_inst_964 (
  .O(mux_o_964),
  .I0(mux_o_959),
  .I1(mux_o_960),
  .S0(dff_q_2)
);
MUX2 mux_inst_965 (
  .O(mux_o_965),
  .I0(mux_o_961),
  .I1(mux_o_962),
  .S0(dff_q_1)
);
MUX2 mux_inst_966 (
  .O(mux_o_966),
  .I0(mux_o_963),
  .I1(mux_o_964),
  .S0(dff_q_1)
);
MUX2 mux_inst_967 (
  .O(dout[7]),
  .I0(mux_o_965),
  .I1(mux_o_966),
  .S0(dff_q_0)
);
MUX2 mux_inst_1027 (
  .O(mux_o_1027),
  .I0(sdpx9b_inst_0_dout[8]),
  .I1(sdpx9b_inst_1_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1028 (
  .O(mux_o_1028),
  .I0(sdpx9b_inst_2_dout[8]),
  .I1(sdpx9b_inst_3_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1029 (
  .O(mux_o_1029),
  .I0(sdpx9b_inst_4_dout[8]),
  .I1(sdpx9b_inst_5_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1030 (
  .O(mux_o_1030),
  .I0(sdpx9b_inst_6_dout[8]),
  .I1(sdpx9b_inst_7_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1031 (
  .O(mux_o_1031),
  .I0(sdpx9b_inst_8_dout[8]),
  .I1(sdpx9b_inst_9_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1032 (
  .O(mux_o_1032),
  .I0(sdpx9b_inst_10_dout[8]),
  .I1(sdpx9b_inst_11_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1033 (
  .O(mux_o_1033),
  .I0(sdpx9b_inst_12_dout[8]),
  .I1(sdpx9b_inst_13_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1034 (
  .O(mux_o_1034),
  .I0(sdpx9b_inst_14_dout[8]),
  .I1(sdpx9b_inst_15_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1035 (
  .O(mux_o_1035),
  .I0(sdpx9b_inst_16_dout[8]),
  .I1(sdpx9b_inst_17_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1036 (
  .O(mux_o_1036),
  .I0(sdpx9b_inst_18_dout[8]),
  .I1(sdpx9b_inst_19_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1037 (
  .O(mux_o_1037),
  .I0(sdpx9b_inst_20_dout[8]),
  .I1(sdpx9b_inst_21_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1038 (
  .O(mux_o_1038),
  .I0(sdpx9b_inst_22_dout[8]),
  .I1(sdpx9b_inst_23_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1039 (
  .O(mux_o_1039),
  .I0(sdpx9b_inst_24_dout[8]),
  .I1(sdpx9b_inst_25_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1040 (
  .O(mux_o_1040),
  .I0(sdpx9b_inst_26_dout[8]),
  .I1(sdpx9b_inst_27_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1041 (
  .O(mux_o_1041),
  .I0(sdpx9b_inst_28_dout[8]),
  .I1(sdpx9b_inst_29_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1042 (
  .O(mux_o_1042),
  .I0(sdpx9b_inst_30_dout[8]),
  .I1(sdpx9b_inst_31_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1043 (
  .O(mux_o_1043),
  .I0(sdpx9b_inst_60_dout[8]),
  .I1(sdpx9b_inst_61_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1044 (
  .O(mux_o_1044),
  .I0(sdpx9b_inst_62_dout[8]),
  .I1(sdpx9b_inst_63_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1045 (
  .O(mux_o_1045),
  .I0(sdpx9b_inst_64_dout[8]),
  .I1(sdpx9b_inst_65_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1046 (
  .O(mux_o_1046),
  .I0(sdpx9b_inst_66_dout[8]),
  .I1(sdpx9b_inst_67_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1047 (
  .O(mux_o_1047),
  .I0(sdpx9b_inst_68_dout[8]),
  .I1(sdpx9b_inst_69_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1048 (
  .O(mux_o_1048),
  .I0(sdpx9b_inst_70_dout[8]),
  .I1(sdpx9b_inst_71_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1049 (
  .O(mux_o_1049),
  .I0(sdpx9b_inst_72_dout[8]),
  .I1(sdpx9b_inst_73_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1050 (
  .O(mux_o_1050),
  .I0(sdpx9b_inst_74_dout[8]),
  .I1(sdpx9b_inst_75_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1051 (
  .O(mux_o_1051),
  .I0(sdpx9b_inst_90_dout[8]),
  .I1(sdpx9b_inst_91_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1052 (
  .O(mux_o_1052),
  .I0(sdpx9b_inst_92_dout[8]),
  .I1(sdpx9b_inst_93_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1053 (
  .O(mux_o_1053),
  .I0(sdpx9b_inst_94_dout[8]),
  .I1(sdpx9b_inst_95_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1054 (
  .O(mux_o_1054),
  .I0(sdpx9b_inst_96_dout[8]),
  .I1(sdpx9b_inst_97_dout[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_1058 (
  .O(mux_o_1058),
  .I0(mux_o_1027),
  .I1(mux_o_1028),
  .S0(dff_q_4)
);
MUX2 mux_inst_1059 (
  .O(mux_o_1059),
  .I0(mux_o_1029),
  .I1(mux_o_1030),
  .S0(dff_q_4)
);
MUX2 mux_inst_1060 (
  .O(mux_o_1060),
  .I0(mux_o_1031),
  .I1(mux_o_1032),
  .S0(dff_q_4)
);
MUX2 mux_inst_1061 (
  .O(mux_o_1061),
  .I0(mux_o_1033),
  .I1(mux_o_1034),
  .S0(dff_q_4)
);
MUX2 mux_inst_1062 (
  .O(mux_o_1062),
  .I0(mux_o_1035),
  .I1(mux_o_1036),
  .S0(dff_q_4)
);
MUX2 mux_inst_1063 (
  .O(mux_o_1063),
  .I0(mux_o_1037),
  .I1(mux_o_1038),
  .S0(dff_q_4)
);
MUX2 mux_inst_1064 (
  .O(mux_o_1064),
  .I0(mux_o_1039),
  .I1(mux_o_1040),
  .S0(dff_q_4)
);
MUX2 mux_inst_1065 (
  .O(mux_o_1065),
  .I0(mux_o_1041),
  .I1(mux_o_1042),
  .S0(dff_q_4)
);
MUX2 mux_inst_1066 (
  .O(mux_o_1066),
  .I0(mux_o_1043),
  .I1(mux_o_1044),
  .S0(dff_q_4)
);
MUX2 mux_inst_1067 (
  .O(mux_o_1067),
  .I0(mux_o_1045),
  .I1(mux_o_1046),
  .S0(dff_q_4)
);
MUX2 mux_inst_1068 (
  .O(mux_o_1068),
  .I0(mux_o_1047),
  .I1(mux_o_1048),
  .S0(dff_q_4)
);
MUX2 mux_inst_1069 (
  .O(mux_o_1069),
  .I0(mux_o_1049),
  .I1(mux_o_1050),
  .S0(dff_q_4)
);
MUX2 mux_inst_1070 (
  .O(mux_o_1070),
  .I0(mux_o_1051),
  .I1(mux_o_1052),
  .S0(dff_q_4)
);
MUX2 mux_inst_1071 (
  .O(mux_o_1071),
  .I0(mux_o_1053),
  .I1(mux_o_1054),
  .S0(dff_q_4)
);
MUX2 mux_inst_1073 (
  .O(mux_o_1073),
  .I0(sdpb_inst_115_dout[8]),
  .I1(sdpb_inst_117_dout[8]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1074 (
  .O(mux_o_1074),
  .I0(mux_o_1058),
  .I1(mux_o_1059),
  .S0(dff_q_3)
);
MUX2 mux_inst_1075 (
  .O(mux_o_1075),
  .I0(mux_o_1060),
  .I1(mux_o_1061),
  .S0(dff_q_3)
);
MUX2 mux_inst_1076 (
  .O(mux_o_1076),
  .I0(mux_o_1062),
  .I1(mux_o_1063),
  .S0(dff_q_3)
);
MUX2 mux_inst_1077 (
  .O(mux_o_1077),
  .I0(mux_o_1064),
  .I1(mux_o_1065),
  .S0(dff_q_3)
);
MUX2 mux_inst_1078 (
  .O(mux_o_1078),
  .I0(mux_o_1066),
  .I1(mux_o_1067),
  .S0(dff_q_3)
);
MUX2 mux_inst_1079 (
  .O(mux_o_1079),
  .I0(mux_o_1068),
  .I1(mux_o_1069),
  .S0(dff_q_3)
);
MUX2 mux_inst_1080 (
  .O(mux_o_1080),
  .I0(mux_o_1070),
  .I1(mux_o_1071),
  .S0(dff_q_3)
);
MUX2 mux_inst_1081 (
  .O(mux_o_1081),
  .I0(sdpb_inst_109_dout[8]),
  .I1(mux_o_1073),
  .S0(dff_q_3)
);
MUX2 mux_inst_1082 (
  .O(mux_o_1082),
  .I0(mux_o_1074),
  .I1(mux_o_1075),
  .S0(dff_q_2)
);
MUX2 mux_inst_1083 (
  .O(mux_o_1083),
  .I0(mux_o_1076),
  .I1(mux_o_1077),
  .S0(dff_q_2)
);
MUX2 mux_inst_1084 (
  .O(mux_o_1084),
  .I0(mux_o_1078),
  .I1(mux_o_1079),
  .S0(dff_q_2)
);
MUX2 mux_inst_1085 (
  .O(mux_o_1085),
  .I0(mux_o_1080),
  .I1(mux_o_1081),
  .S0(dff_q_2)
);
MUX2 mux_inst_1086 (
  .O(mux_o_1086),
  .I0(mux_o_1082),
  .I1(mux_o_1083),
  .S0(dff_q_1)
);
MUX2 mux_inst_1087 (
  .O(mux_o_1087),
  .I0(mux_o_1084),
  .I1(mux_o_1085),
  .S0(dff_q_1)
);
MUX2 mux_inst_1088 (
  .O(dout[8]),
  .I0(mux_o_1086),
  .I1(mux_o_1087),
  .S0(dff_q_0)
);
MUX2 mux_inst_1117 (
  .O(mux_o_1117),
  .I0(sdpb_inst_115_dout[9]),
  .I1(sdpb_inst_117_dout[9]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1125 (
  .O(mux_o_1125),
  .I0(sdpb_inst_109_dout[9]),
  .I1(mux_o_1117),
  .S0(dff_q_3)
);
MUX2 mux_inst_1126 (
  .O(mux_o_1126),
  .I0(sdpb_inst_32_dout[9]),
  .I1(sdpb_inst_33_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1127 (
  .O(mux_o_1127),
  .I0(sdpb_inst_34_dout[9]),
  .I1(sdpb_inst_35_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1128 (
  .O(mux_o_1128),
  .I0(sdpb_inst_76_dout[9]),
  .I1(sdpb_inst_77_dout[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1129 (
  .O(mux_o_1129),
  .I0(sdpb_inst_98_dout[9]),
  .I1(mux_o_1125),
  .S0(dff_q_2)
);
MUX2 mux_inst_1130 (
  .O(mux_o_1130),
  .I0(mux_o_1126),
  .I1(mux_o_1127),
  .S0(dff_q_1)
);
MUX2 mux_inst_1131 (
  .O(mux_o_1131),
  .I0(mux_o_1128),
  .I1(mux_o_1129),
  .S0(dff_q_1)
);
MUX2 mux_inst_1132 (
  .O(dout[9]),
  .I0(mux_o_1130),
  .I1(mux_o_1131),
  .S0(dff_q_0)
);
MUX2 mux_inst_1161 (
  .O(mux_o_1161),
  .I0(sdpb_inst_115_dout[10]),
  .I1(sdpb_inst_117_dout[10]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1169 (
  .O(mux_o_1169),
  .I0(sdpb_inst_110_dout[10]),
  .I1(mux_o_1161),
  .S0(dff_q_3)
);
MUX2 mux_inst_1170 (
  .O(mux_o_1170),
  .I0(sdpb_inst_36_dout[10]),
  .I1(sdpb_inst_37_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1171 (
  .O(mux_o_1171),
  .I0(sdpb_inst_38_dout[10]),
  .I1(sdpb_inst_39_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1172 (
  .O(mux_o_1172),
  .I0(sdpb_inst_78_dout[10]),
  .I1(sdpb_inst_79_dout[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1173 (
  .O(mux_o_1173),
  .I0(sdpb_inst_99_dout[10]),
  .I1(mux_o_1169),
  .S0(dff_q_2)
);
MUX2 mux_inst_1174 (
  .O(mux_o_1174),
  .I0(mux_o_1170),
  .I1(mux_o_1171),
  .S0(dff_q_1)
);
MUX2 mux_inst_1175 (
  .O(mux_o_1175),
  .I0(mux_o_1172),
  .I1(mux_o_1173),
  .S0(dff_q_1)
);
MUX2 mux_inst_1176 (
  .O(dout[10]),
  .I0(mux_o_1174),
  .I1(mux_o_1175),
  .S0(dff_q_0)
);
MUX2 mux_inst_1205 (
  .O(mux_o_1205),
  .I0(sdpb_inst_115_dout[11]),
  .I1(sdpb_inst_117_dout[11]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1213 (
  .O(mux_o_1213),
  .I0(sdpb_inst_110_dout[11]),
  .I1(mux_o_1205),
  .S0(dff_q_3)
);
MUX2 mux_inst_1214 (
  .O(mux_o_1214),
  .I0(sdpb_inst_40_dout[11]),
  .I1(sdpb_inst_41_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1215 (
  .O(mux_o_1215),
  .I0(sdpb_inst_42_dout[11]),
  .I1(sdpb_inst_43_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1216 (
  .O(mux_o_1216),
  .I0(sdpb_inst_80_dout[11]),
  .I1(sdpb_inst_81_dout[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1217 (
  .O(mux_o_1217),
  .I0(sdpb_inst_100_dout[11]),
  .I1(mux_o_1213),
  .S0(dff_q_2)
);
MUX2 mux_inst_1218 (
  .O(mux_o_1218),
  .I0(mux_o_1214),
  .I1(mux_o_1215),
  .S0(dff_q_1)
);
MUX2 mux_inst_1219 (
  .O(mux_o_1219),
  .I0(mux_o_1216),
  .I1(mux_o_1217),
  .S0(dff_q_1)
);
MUX2 mux_inst_1220 (
  .O(dout[11]),
  .I0(mux_o_1218),
  .I1(mux_o_1219),
  .S0(dff_q_0)
);
MUX2 mux_inst_1249 (
  .O(mux_o_1249),
  .I0(sdpb_inst_116_dout[12]),
  .I1(sdpb_inst_117_dout[12]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1257 (
  .O(mux_o_1257),
  .I0(sdpb_inst_111_dout[12]),
  .I1(mux_o_1249),
  .S0(dff_q_3)
);
MUX2 mux_inst_1258 (
  .O(mux_o_1258),
  .I0(sdpb_inst_44_dout[12]),
  .I1(sdpb_inst_45_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1259 (
  .O(mux_o_1259),
  .I0(sdpb_inst_46_dout[12]),
  .I1(sdpb_inst_47_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1260 (
  .O(mux_o_1260),
  .I0(sdpb_inst_82_dout[12]),
  .I1(sdpb_inst_83_dout[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1261 (
  .O(mux_o_1261),
  .I0(sdpb_inst_101_dout[12]),
  .I1(mux_o_1257),
  .S0(dff_q_2)
);
MUX2 mux_inst_1262 (
  .O(mux_o_1262),
  .I0(mux_o_1258),
  .I1(mux_o_1259),
  .S0(dff_q_1)
);
MUX2 mux_inst_1263 (
  .O(mux_o_1263),
  .I0(mux_o_1260),
  .I1(mux_o_1261),
  .S0(dff_q_1)
);
MUX2 mux_inst_1264 (
  .O(dout[12]),
  .I0(mux_o_1262),
  .I1(mux_o_1263),
  .S0(dff_q_0)
);
MUX2 mux_inst_1293 (
  .O(mux_o_1293),
  .I0(sdpb_inst_116_dout[13]),
  .I1(sdpb_inst_117_dout[13]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1301 (
  .O(mux_o_1301),
  .I0(sdpb_inst_111_dout[13]),
  .I1(mux_o_1293),
  .S0(dff_q_3)
);
MUX2 mux_inst_1302 (
  .O(mux_o_1302),
  .I0(sdpb_inst_48_dout[13]),
  .I1(sdpb_inst_49_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1303 (
  .O(mux_o_1303),
  .I0(sdpb_inst_50_dout[13]),
  .I1(sdpb_inst_51_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1304 (
  .O(mux_o_1304),
  .I0(sdpb_inst_84_dout[13]),
  .I1(sdpb_inst_85_dout[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1305 (
  .O(mux_o_1305),
  .I0(sdpb_inst_102_dout[13]),
  .I1(mux_o_1301),
  .S0(dff_q_2)
);
MUX2 mux_inst_1306 (
  .O(mux_o_1306),
  .I0(mux_o_1302),
  .I1(mux_o_1303),
  .S0(dff_q_1)
);
MUX2 mux_inst_1307 (
  .O(mux_o_1307),
  .I0(mux_o_1304),
  .I1(mux_o_1305),
  .S0(dff_q_1)
);
MUX2 mux_inst_1308 (
  .O(dout[13]),
  .I0(mux_o_1306),
  .I1(mux_o_1307),
  .S0(dff_q_0)
);
MUX2 mux_inst_1337 (
  .O(mux_o_1337),
  .I0(sdpb_inst_116_dout[14]),
  .I1(sdpb_inst_117_dout[14]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1345 (
  .O(mux_o_1345),
  .I0(sdpb_inst_112_dout[14]),
  .I1(mux_o_1337),
  .S0(dff_q_3)
);
MUX2 mux_inst_1346 (
  .O(mux_o_1346),
  .I0(sdpb_inst_52_dout[14]),
  .I1(sdpb_inst_53_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1347 (
  .O(mux_o_1347),
  .I0(sdpb_inst_54_dout[14]),
  .I1(sdpb_inst_55_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1348 (
  .O(mux_o_1348),
  .I0(sdpb_inst_86_dout[14]),
  .I1(sdpb_inst_87_dout[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1349 (
  .O(mux_o_1349),
  .I0(sdpb_inst_103_dout[14]),
  .I1(mux_o_1345),
  .S0(dff_q_2)
);
MUX2 mux_inst_1350 (
  .O(mux_o_1350),
  .I0(mux_o_1346),
  .I1(mux_o_1347),
  .S0(dff_q_1)
);
MUX2 mux_inst_1351 (
  .O(mux_o_1351),
  .I0(mux_o_1348),
  .I1(mux_o_1349),
  .S0(dff_q_1)
);
MUX2 mux_inst_1352 (
  .O(dout[14]),
  .I0(mux_o_1350),
  .I1(mux_o_1351),
  .S0(dff_q_0)
);
MUX2 mux_inst_1381 (
  .O(mux_o_1381),
  .I0(sdpb_inst_116_dout[15]),
  .I1(sdpb_inst_117_dout[15]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1389 (
  .O(mux_o_1389),
  .I0(sdpb_inst_112_dout[15]),
  .I1(mux_o_1381),
  .S0(dff_q_3)
);
MUX2 mux_inst_1390 (
  .O(mux_o_1390),
  .I0(sdpb_inst_56_dout[15]),
  .I1(sdpb_inst_57_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1391 (
  .O(mux_o_1391),
  .I0(sdpb_inst_58_dout[15]),
  .I1(sdpb_inst_59_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1392 (
  .O(mux_o_1392),
  .I0(sdpb_inst_88_dout[15]),
  .I1(sdpb_inst_89_dout[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1393 (
  .O(mux_o_1393),
  .I0(sdpb_inst_104_dout[15]),
  .I1(mux_o_1389),
  .S0(dff_q_2)
);
MUX2 mux_inst_1394 (
  .O(mux_o_1394),
  .I0(mux_o_1390),
  .I1(mux_o_1391),
  .S0(dff_q_1)
);
MUX2 mux_inst_1395 (
  .O(mux_o_1395),
  .I0(mux_o_1392),
  .I1(mux_o_1393),
  .S0(dff_q_1)
);
MUX2 mux_inst_1396 (
  .O(dout[15]),
  .I0(mux_o_1394),
  .I1(mux_o_1395),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB
